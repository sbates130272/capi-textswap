`default_nettype none
//------------------------------------------------------------------
//-- This module implements a 128-bit external LFSR that advances --
//-- 512 states per clock. The polynomial for this LFSR is given  --
//-- as: p(x) = x^128 + x^126 + x^101 + x^99 + 1                  --
//--                                                              --
//-- Saeed Fouladi Fard, PhD, PMC-Sierra                          --
//------------------------------------------------------------------

module lfsr
 (
   input  wire           clk      ,   // clock, rising edge
   input  wire           reset    ,   // reset, sync, active high. At reset the LFSR is set to all ones
   input  wire [128-1:0] i_seed   ,   // LFSR seed, picked when init=1
   input  wire           i_init   ,   // When high, the LFSR will be seeded with seed. i_init overrides i_advance
   input  wire           i_advance,   // When high, state of the LFSR advances by 512 steps
   output wire  [512-1:0] o_lfsr      // State of the LFSR
 );

  // Internal signals:
  reg     [128-1:0] lfsr;
  initial lfsr = {(512){1'b1}};
  integer           i;


  // XOR-tree for the LFSR

  assign  o_lfsr[ 0] = lfsr[98]^lfsr[100]^lfsr[125]^lfsr[127];
  assign  o_lfsr[ 1] = lfsr[97]^lfsr[99]^lfsr[124]^lfsr[126];
  assign  o_lfsr[ 2] = lfsr[96]^lfsr[98]^lfsr[123]^lfsr[125];
  assign  o_lfsr[ 3] = lfsr[95]^lfsr[97]^lfsr[122]^lfsr[124];
  assign  o_lfsr[ 4] = lfsr[94]^lfsr[96]^lfsr[121]^lfsr[123];
  assign  o_lfsr[ 5] = lfsr[93]^lfsr[95]^lfsr[120]^lfsr[122];
  assign  o_lfsr[ 6] = lfsr[92]^lfsr[94]^lfsr[119]^lfsr[121];
  assign  o_lfsr[ 7] = lfsr[91]^lfsr[93]^lfsr[118]^lfsr[120];
  assign  o_lfsr[ 8] = lfsr[90]^lfsr[92]^lfsr[117]^lfsr[119];
  assign  o_lfsr[ 9] = lfsr[89]^lfsr[91]^lfsr[116]^lfsr[118];
  assign  o_lfsr[10] = lfsr[88]^lfsr[90]^lfsr[115]^lfsr[117];
  assign  o_lfsr[11] = lfsr[87]^lfsr[89]^lfsr[114]^lfsr[116];
  assign  o_lfsr[12] = lfsr[86]^lfsr[88]^lfsr[113]^lfsr[115];
  assign  o_lfsr[13] = lfsr[85]^lfsr[87]^lfsr[112]^lfsr[114];
  assign  o_lfsr[14] = lfsr[84]^lfsr[86]^lfsr[111]^lfsr[113];
  assign  o_lfsr[15] = lfsr[83]^lfsr[85]^lfsr[110]^lfsr[112];
  assign  o_lfsr[16] = lfsr[82]^lfsr[84]^lfsr[109]^lfsr[111];
  assign  o_lfsr[17] = lfsr[81]^lfsr[83]^lfsr[108]^lfsr[110];
  assign  o_lfsr[18] = lfsr[80]^lfsr[82]^lfsr[107]^lfsr[109];
  assign  o_lfsr[19] = lfsr[79]^lfsr[81]^lfsr[106]^lfsr[108];
  assign  o_lfsr[20] = lfsr[78]^lfsr[80]^lfsr[105]^lfsr[107];
  assign  o_lfsr[21] = lfsr[77]^lfsr[79]^lfsr[104]^lfsr[106];
  assign  o_lfsr[22] = lfsr[76]^lfsr[78]^lfsr[103]^lfsr[105];
  assign  o_lfsr[23] = lfsr[75]^lfsr[77]^lfsr[102]^lfsr[104];
  assign  o_lfsr[24] = lfsr[74]^lfsr[76]^lfsr[101]^lfsr[103];
  assign  o_lfsr[25] = lfsr[73]^lfsr[75]^lfsr[100]^lfsr[102];
  assign  o_lfsr[26] = lfsr[72]^lfsr[74]^lfsr[99]^lfsr[101];
  assign  o_lfsr[27] = lfsr[71]^lfsr[73]^lfsr[98]^lfsr[100];
  assign  o_lfsr[28] = lfsr[70]^lfsr[72]^lfsr[97]^lfsr[99];
  assign  o_lfsr[29] = lfsr[69]^lfsr[71]^lfsr[96]^lfsr[98];
  assign  o_lfsr[30] = lfsr[68]^lfsr[70]^lfsr[95]^lfsr[97];
  assign  o_lfsr[31] = lfsr[67]^lfsr[69]^lfsr[94]^lfsr[96];
  assign  o_lfsr[32] = lfsr[66]^lfsr[68]^lfsr[93]^lfsr[95];
  assign  o_lfsr[33] = lfsr[65]^lfsr[67]^lfsr[92]^lfsr[94];
  assign  o_lfsr[34] = lfsr[64]^lfsr[66]^lfsr[91]^lfsr[93];
  assign  o_lfsr[35] = lfsr[63]^lfsr[65]^lfsr[90]^lfsr[92];
  assign  o_lfsr[36] = lfsr[62]^lfsr[64]^lfsr[89]^lfsr[91];
  assign  o_lfsr[37] = lfsr[61]^lfsr[63]^lfsr[88]^lfsr[90];
  assign  o_lfsr[38] = lfsr[60]^lfsr[62]^lfsr[87]^lfsr[89];
  assign  o_lfsr[39] = lfsr[59]^lfsr[61]^lfsr[86]^lfsr[88];
  assign  o_lfsr[40] = lfsr[58]^lfsr[60]^lfsr[85]^lfsr[87];
  assign  o_lfsr[41] = lfsr[57]^lfsr[59]^lfsr[84]^lfsr[86];
  assign  o_lfsr[42] = lfsr[56]^lfsr[58]^lfsr[83]^lfsr[85];
  assign  o_lfsr[43] = lfsr[55]^lfsr[57]^lfsr[82]^lfsr[84];
  assign  o_lfsr[44] = lfsr[54]^lfsr[56]^lfsr[81]^lfsr[83];
  assign  o_lfsr[45] = lfsr[53]^lfsr[55]^lfsr[80]^lfsr[82];
  assign  o_lfsr[46] = lfsr[52]^lfsr[54]^lfsr[79]^lfsr[81];
  assign  o_lfsr[47] = lfsr[51]^lfsr[53]^lfsr[78]^lfsr[80];
  assign  o_lfsr[48] = lfsr[50]^lfsr[52]^lfsr[77]^lfsr[79];
  assign  o_lfsr[49] = lfsr[49]^lfsr[51]^lfsr[76]^lfsr[78];
  assign  o_lfsr[50] = lfsr[48]^lfsr[50]^lfsr[75]^lfsr[77];
  assign  o_lfsr[51] = lfsr[47]^lfsr[49]^lfsr[74]^lfsr[76];
  assign  o_lfsr[52] = lfsr[46]^lfsr[48]^lfsr[73]^lfsr[75];
  assign  o_lfsr[53] = lfsr[45]^lfsr[47]^lfsr[72]^lfsr[74];
  assign  o_lfsr[54] = lfsr[44]^lfsr[46]^lfsr[71]^lfsr[73];
  assign  o_lfsr[55] = lfsr[43]^lfsr[45]^lfsr[70]^lfsr[72];
  assign  o_lfsr[56] = lfsr[42]^lfsr[44]^lfsr[69]^lfsr[71];
  assign  o_lfsr[57] = lfsr[41]^lfsr[43]^lfsr[68]^lfsr[70];
  assign  o_lfsr[58] = lfsr[40]^lfsr[42]^lfsr[67]^lfsr[69];
  assign  o_lfsr[59] = lfsr[39]^lfsr[41]^lfsr[66]^lfsr[68];
  assign  o_lfsr[60] = lfsr[38]^lfsr[40]^lfsr[65]^lfsr[67];
  assign  o_lfsr[61] = lfsr[37]^lfsr[39]^lfsr[64]^lfsr[66];
  assign  o_lfsr[62] = lfsr[36]^lfsr[38]^lfsr[63]^lfsr[65];
  assign  o_lfsr[63] = lfsr[35]^lfsr[37]^lfsr[62]^lfsr[64];
  assign  o_lfsr[64] = lfsr[34]^lfsr[36]^lfsr[61]^lfsr[63];
  assign  o_lfsr[65] = lfsr[33]^lfsr[35]^lfsr[60]^lfsr[62];
  assign  o_lfsr[66] = lfsr[32]^lfsr[34]^lfsr[59]^lfsr[61];
  assign  o_lfsr[67] = lfsr[31]^lfsr[33]^lfsr[58]^lfsr[60];
  assign  o_lfsr[68] = lfsr[30]^lfsr[32]^lfsr[57]^lfsr[59];
  assign  o_lfsr[69] = lfsr[29]^lfsr[31]^lfsr[56]^lfsr[58];
  assign  o_lfsr[70] = lfsr[28]^lfsr[30]^lfsr[55]^lfsr[57];
  assign  o_lfsr[71] = lfsr[27]^lfsr[29]^lfsr[54]^lfsr[56];
  assign  o_lfsr[72] = lfsr[26]^lfsr[28]^lfsr[53]^lfsr[55];
  assign  o_lfsr[73] = lfsr[25]^lfsr[27]^lfsr[52]^lfsr[54];
  assign  o_lfsr[74] = lfsr[24]^lfsr[26]^lfsr[51]^lfsr[53];
  assign  o_lfsr[75] = lfsr[23]^lfsr[25]^lfsr[50]^lfsr[52];
  assign  o_lfsr[76] = lfsr[22]^lfsr[24]^lfsr[49]^lfsr[51];
  assign  o_lfsr[77] = lfsr[21]^lfsr[23]^lfsr[48]^lfsr[50];
  assign  o_lfsr[78] = lfsr[20]^lfsr[22]^lfsr[47]^lfsr[49];
  assign  o_lfsr[79] = lfsr[19]^lfsr[21]^lfsr[46]^lfsr[48];
  assign  o_lfsr[80] = lfsr[18]^lfsr[20]^lfsr[45]^lfsr[47];
  assign  o_lfsr[81] = lfsr[17]^lfsr[19]^lfsr[44]^lfsr[46];
  assign  o_lfsr[82] = lfsr[16]^lfsr[18]^lfsr[43]^lfsr[45];
  assign  o_lfsr[83] = lfsr[15]^lfsr[17]^lfsr[42]^lfsr[44];
  assign  o_lfsr[84] = lfsr[14]^lfsr[16]^lfsr[41]^lfsr[43];
  assign  o_lfsr[85] = lfsr[13]^lfsr[15]^lfsr[40]^lfsr[42];
  assign  o_lfsr[86] = lfsr[12]^lfsr[14]^lfsr[39]^lfsr[41];
  assign  o_lfsr[87] = lfsr[11]^lfsr[13]^lfsr[38]^lfsr[40];
  assign  o_lfsr[88] = lfsr[10]^lfsr[12]^lfsr[37]^lfsr[39];
  assign  o_lfsr[89] = lfsr[ 9]^lfsr[11]^lfsr[36]^lfsr[38];
  assign  o_lfsr[90] = lfsr[ 8]^lfsr[10]^lfsr[35]^lfsr[37];
  assign  o_lfsr[91] = lfsr[ 7]^lfsr[ 9]^lfsr[34]^lfsr[36];
  assign  o_lfsr[92] = lfsr[ 6]^lfsr[ 8]^lfsr[33]^lfsr[35];
  assign  o_lfsr[93] = lfsr[ 5]^lfsr[ 7]^lfsr[32]^lfsr[34];
  assign  o_lfsr[94] = lfsr[ 4]^lfsr[ 6]^lfsr[31]^lfsr[33];
  assign  o_lfsr[95] = lfsr[ 3]^lfsr[ 5]^lfsr[30]^lfsr[32];
  assign  o_lfsr[96] = lfsr[ 2]^lfsr[ 4]^lfsr[29]^lfsr[31];
  assign  o_lfsr[97] = lfsr[ 1]^lfsr[ 3]^lfsr[28]^lfsr[30];
  assign  o_lfsr[98] = lfsr[ 0]^lfsr[ 2]^lfsr[27]^lfsr[29];
  assign  o_lfsr[99] = lfsr[ 1]^lfsr[26]^lfsr[28]^lfsr[98]^lfsr[100]^lfsr[125]^lfsr[127];
  assign  o_lfsr[100] = lfsr[ 0]^lfsr[25]^lfsr[27]^lfsr[97]^lfsr[99]^lfsr[124]^lfsr[126];
  assign  o_lfsr[101] = lfsr[24]^lfsr[26]^lfsr[96]^lfsr[100]^lfsr[123]^lfsr[127];
  assign  o_lfsr[102] = lfsr[23]^lfsr[25]^lfsr[95]^lfsr[99]^lfsr[122]^lfsr[126];
  assign  o_lfsr[103] = lfsr[22]^lfsr[24]^lfsr[94]^lfsr[98]^lfsr[121]^lfsr[125];
  assign  o_lfsr[104] = lfsr[21]^lfsr[23]^lfsr[93]^lfsr[97]^lfsr[120]^lfsr[124];
  assign  o_lfsr[105] = lfsr[20]^lfsr[22]^lfsr[92]^lfsr[96]^lfsr[119]^lfsr[123];
  assign  o_lfsr[106] = lfsr[19]^lfsr[21]^lfsr[91]^lfsr[95]^lfsr[118]^lfsr[122];
  assign  o_lfsr[107] = lfsr[18]^lfsr[20]^lfsr[90]^lfsr[94]^lfsr[117]^lfsr[121];
  assign  o_lfsr[108] = lfsr[17]^lfsr[19]^lfsr[89]^lfsr[93]^lfsr[116]^lfsr[120];
  assign  o_lfsr[109] = lfsr[16]^lfsr[18]^lfsr[88]^lfsr[92]^lfsr[115]^lfsr[119];
  assign  o_lfsr[110] = lfsr[15]^lfsr[17]^lfsr[87]^lfsr[91]^lfsr[114]^lfsr[118];
  assign  o_lfsr[111] = lfsr[14]^lfsr[16]^lfsr[86]^lfsr[90]^lfsr[113]^lfsr[117];
  assign  o_lfsr[112] = lfsr[13]^lfsr[15]^lfsr[85]^lfsr[89]^lfsr[112]^lfsr[116];
  assign  o_lfsr[113] = lfsr[12]^lfsr[14]^lfsr[84]^lfsr[88]^lfsr[111]^lfsr[115];
  assign  o_lfsr[114] = lfsr[11]^lfsr[13]^lfsr[83]^lfsr[87]^lfsr[110]^lfsr[114];
  assign  o_lfsr[115] = lfsr[10]^lfsr[12]^lfsr[82]^lfsr[86]^lfsr[109]^lfsr[113];
  assign  o_lfsr[116] = lfsr[ 9]^lfsr[11]^lfsr[81]^lfsr[85]^lfsr[108]^lfsr[112];
  assign  o_lfsr[117] = lfsr[ 8]^lfsr[10]^lfsr[80]^lfsr[84]^lfsr[107]^lfsr[111];
  assign  o_lfsr[118] = lfsr[ 7]^lfsr[ 9]^lfsr[79]^lfsr[83]^lfsr[106]^lfsr[110];
  assign  o_lfsr[119] = lfsr[ 6]^lfsr[ 8]^lfsr[78]^lfsr[82]^lfsr[105]^lfsr[109];
  assign  o_lfsr[120] = lfsr[ 5]^lfsr[ 7]^lfsr[77]^lfsr[81]^lfsr[104]^lfsr[108];
  assign  o_lfsr[121] = lfsr[ 4]^lfsr[ 6]^lfsr[76]^lfsr[80]^lfsr[103]^lfsr[107];
  assign  o_lfsr[122] = lfsr[ 3]^lfsr[ 5]^lfsr[75]^lfsr[79]^lfsr[102]^lfsr[106];
  assign  o_lfsr[123] = lfsr[ 2]^lfsr[ 4]^lfsr[74]^lfsr[78]^lfsr[101]^lfsr[105];
  assign  o_lfsr[124] = lfsr[ 1]^lfsr[ 3]^lfsr[73]^lfsr[77]^lfsr[100]^lfsr[104];
  assign  o_lfsr[125] = lfsr[ 0]^lfsr[ 2]^lfsr[72]^lfsr[76]^lfsr[99]^lfsr[103];
  assign  o_lfsr[126] = lfsr[ 1]^lfsr[71]^lfsr[75]^lfsr[100]^lfsr[102]^lfsr[125]^lfsr[127];
  assign  o_lfsr[127] = lfsr[ 0]^lfsr[70]^lfsr[74]^lfsr[99]^lfsr[101]^lfsr[124]^lfsr[126];
  assign  o_lfsr[128] = lfsr[69]^lfsr[73]^lfsr[123]^lfsr[127];
  assign  o_lfsr[129] = lfsr[68]^lfsr[72]^lfsr[122]^lfsr[126];
  assign  o_lfsr[130] = lfsr[67]^lfsr[71]^lfsr[121]^lfsr[125];
  assign  o_lfsr[131] = lfsr[66]^lfsr[70]^lfsr[120]^lfsr[124];
  assign  o_lfsr[132] = lfsr[65]^lfsr[69]^lfsr[119]^lfsr[123];
  assign  o_lfsr[133] = lfsr[64]^lfsr[68]^lfsr[118]^lfsr[122];
  assign  o_lfsr[134] = lfsr[63]^lfsr[67]^lfsr[117]^lfsr[121];
  assign  o_lfsr[135] = lfsr[62]^lfsr[66]^lfsr[116]^lfsr[120];
  assign  o_lfsr[136] = lfsr[61]^lfsr[65]^lfsr[115]^lfsr[119];
  assign  o_lfsr[137] = lfsr[60]^lfsr[64]^lfsr[114]^lfsr[118];
  assign  o_lfsr[138] = lfsr[59]^lfsr[63]^lfsr[113]^lfsr[117];
  assign  o_lfsr[139] = lfsr[58]^lfsr[62]^lfsr[112]^lfsr[116];
  assign  o_lfsr[140] = lfsr[57]^lfsr[61]^lfsr[111]^lfsr[115];
  assign  o_lfsr[141] = lfsr[56]^lfsr[60]^lfsr[110]^lfsr[114];
  assign  o_lfsr[142] = lfsr[55]^lfsr[59]^lfsr[109]^lfsr[113];
  assign  o_lfsr[143] = lfsr[54]^lfsr[58]^lfsr[108]^lfsr[112];
  assign  o_lfsr[144] = lfsr[53]^lfsr[57]^lfsr[107]^lfsr[111];
  assign  o_lfsr[145] = lfsr[52]^lfsr[56]^lfsr[106]^lfsr[110];
  assign  o_lfsr[146] = lfsr[51]^lfsr[55]^lfsr[105]^lfsr[109];
  assign  o_lfsr[147] = lfsr[50]^lfsr[54]^lfsr[104]^lfsr[108];
  assign  o_lfsr[148] = lfsr[49]^lfsr[53]^lfsr[103]^lfsr[107];
  assign  o_lfsr[149] = lfsr[48]^lfsr[52]^lfsr[102]^lfsr[106];
  assign  o_lfsr[150] = lfsr[47]^lfsr[51]^lfsr[101]^lfsr[105];
  assign  o_lfsr[151] = lfsr[46]^lfsr[50]^lfsr[100]^lfsr[104];
  assign  o_lfsr[152] = lfsr[45]^lfsr[49]^lfsr[99]^lfsr[103];
  assign  o_lfsr[153] = lfsr[44]^lfsr[48]^lfsr[98]^lfsr[102];
  assign  o_lfsr[154] = lfsr[43]^lfsr[47]^lfsr[97]^lfsr[101];
  assign  o_lfsr[155] = lfsr[42]^lfsr[46]^lfsr[96]^lfsr[100];
  assign  o_lfsr[156] = lfsr[41]^lfsr[45]^lfsr[95]^lfsr[99];
  assign  o_lfsr[157] = lfsr[40]^lfsr[44]^lfsr[94]^lfsr[98];
  assign  o_lfsr[158] = lfsr[39]^lfsr[43]^lfsr[93]^lfsr[97];
  assign  o_lfsr[159] = lfsr[38]^lfsr[42]^lfsr[92]^lfsr[96];
  assign  o_lfsr[160] = lfsr[37]^lfsr[41]^lfsr[91]^lfsr[95];
  assign  o_lfsr[161] = lfsr[36]^lfsr[40]^lfsr[90]^lfsr[94];
  assign  o_lfsr[162] = lfsr[35]^lfsr[39]^lfsr[89]^lfsr[93];
  assign  o_lfsr[163] = lfsr[34]^lfsr[38]^lfsr[88]^lfsr[92];
  assign  o_lfsr[164] = lfsr[33]^lfsr[37]^lfsr[87]^lfsr[91];
  assign  o_lfsr[165] = lfsr[32]^lfsr[36]^lfsr[86]^lfsr[90];
  assign  o_lfsr[166] = lfsr[31]^lfsr[35]^lfsr[85]^lfsr[89];
  assign  o_lfsr[167] = lfsr[30]^lfsr[34]^lfsr[84]^lfsr[88];
  assign  o_lfsr[168] = lfsr[29]^lfsr[33]^lfsr[83]^lfsr[87];
  assign  o_lfsr[169] = lfsr[28]^lfsr[32]^lfsr[82]^lfsr[86];
  assign  o_lfsr[170] = lfsr[27]^lfsr[31]^lfsr[81]^lfsr[85];
  assign  o_lfsr[171] = lfsr[26]^lfsr[30]^lfsr[80]^lfsr[84];
  assign  o_lfsr[172] = lfsr[25]^lfsr[29]^lfsr[79]^lfsr[83];
  assign  o_lfsr[173] = lfsr[24]^lfsr[28]^lfsr[78]^lfsr[82];
  assign  o_lfsr[174] = lfsr[23]^lfsr[27]^lfsr[77]^lfsr[81];
  assign  o_lfsr[175] = lfsr[22]^lfsr[26]^lfsr[76]^lfsr[80];
  assign  o_lfsr[176] = lfsr[21]^lfsr[25]^lfsr[75]^lfsr[79];
  assign  o_lfsr[177] = lfsr[20]^lfsr[24]^lfsr[74]^lfsr[78];
  assign  o_lfsr[178] = lfsr[19]^lfsr[23]^lfsr[73]^lfsr[77];
  assign  o_lfsr[179] = lfsr[18]^lfsr[22]^lfsr[72]^lfsr[76];
  assign  o_lfsr[180] = lfsr[17]^lfsr[21]^lfsr[71]^lfsr[75];
  assign  o_lfsr[181] = lfsr[16]^lfsr[20]^lfsr[70]^lfsr[74];
  assign  o_lfsr[182] = lfsr[15]^lfsr[19]^lfsr[69]^lfsr[73];
  assign  o_lfsr[183] = lfsr[14]^lfsr[18]^lfsr[68]^lfsr[72];
  assign  o_lfsr[184] = lfsr[13]^lfsr[17]^lfsr[67]^lfsr[71];
  assign  o_lfsr[185] = lfsr[12]^lfsr[16]^lfsr[66]^lfsr[70];
  assign  o_lfsr[186] = lfsr[11]^lfsr[15]^lfsr[65]^lfsr[69];
  assign  o_lfsr[187] = lfsr[10]^lfsr[14]^lfsr[64]^lfsr[68];
  assign  o_lfsr[188] = lfsr[ 9]^lfsr[13]^lfsr[63]^lfsr[67];
  assign  o_lfsr[189] = lfsr[ 8]^lfsr[12]^lfsr[62]^lfsr[66];
  assign  o_lfsr[190] = lfsr[ 7]^lfsr[11]^lfsr[61]^lfsr[65];
  assign  o_lfsr[191] = lfsr[ 6]^lfsr[10]^lfsr[60]^lfsr[64];
  assign  o_lfsr[192] = lfsr[ 5]^lfsr[ 9]^lfsr[59]^lfsr[63];
  assign  o_lfsr[193] = lfsr[ 4]^lfsr[ 8]^lfsr[58]^lfsr[62];
  assign  o_lfsr[194] = lfsr[ 3]^lfsr[ 7]^lfsr[57]^lfsr[61];
  assign  o_lfsr[195] = lfsr[ 2]^lfsr[ 6]^lfsr[56]^lfsr[60];
  assign  o_lfsr[196] = lfsr[ 1]^lfsr[ 5]^lfsr[55]^lfsr[59];
  assign  o_lfsr[197] = lfsr[ 0]^lfsr[ 4]^lfsr[54]^lfsr[58];
  assign  o_lfsr[198] = lfsr[ 3]^lfsr[53]^lfsr[57]^lfsr[98]^lfsr[100]^lfsr[125]^lfsr[127];
  assign  o_lfsr[199] = lfsr[ 2]^lfsr[52]^lfsr[56]^lfsr[97]^lfsr[99]^lfsr[124]^lfsr[126];
  assign  o_lfsr[200] = lfsr[ 1]^lfsr[51]^lfsr[55]^lfsr[96]^lfsr[98]^lfsr[123]^lfsr[125];
  assign  o_lfsr[201] = lfsr[ 0]^lfsr[50]^lfsr[54]^lfsr[95]^lfsr[97]^lfsr[122]^lfsr[124];
  assign  o_lfsr[202] = lfsr[49]^lfsr[53]^lfsr[94]^lfsr[96]^lfsr[98]^lfsr[100]^lfsr[121]^lfsr[123]^lfsr[125]^lfsr[127];
  assign  o_lfsr[203] = lfsr[48]^lfsr[52]^lfsr[93]^lfsr[95]^lfsr[97]^lfsr[99]^lfsr[120]^lfsr[122]^lfsr[124]^lfsr[126];
  assign  o_lfsr[204] = lfsr[47]^lfsr[51]^lfsr[92]^lfsr[94]^lfsr[96]^lfsr[98]^lfsr[119]^lfsr[121]^lfsr[123]^lfsr[125];
  assign  o_lfsr[205] = lfsr[46]^lfsr[50]^lfsr[91]^lfsr[93]^lfsr[95]^lfsr[97]^lfsr[118]^lfsr[120]^lfsr[122]^lfsr[124];
  assign  o_lfsr[206] = lfsr[45]^lfsr[49]^lfsr[90]^lfsr[92]^lfsr[94]^lfsr[96]^lfsr[117]^lfsr[119]^lfsr[121]^lfsr[123];
  assign  o_lfsr[207] = lfsr[44]^lfsr[48]^lfsr[89]^lfsr[91]^lfsr[93]^lfsr[95]^lfsr[116]^lfsr[118]^lfsr[120]^lfsr[122];
  assign  o_lfsr[208] = lfsr[43]^lfsr[47]^lfsr[88]^lfsr[90]^lfsr[92]^lfsr[94]^lfsr[115]^lfsr[117]^lfsr[119]^lfsr[121];
  assign  o_lfsr[209] = lfsr[42]^lfsr[46]^lfsr[87]^lfsr[89]^lfsr[91]^lfsr[93]^lfsr[114]^lfsr[116]^lfsr[118]^lfsr[120];
  assign  o_lfsr[210] = lfsr[41]^lfsr[45]^lfsr[86]^lfsr[88]^lfsr[90]^lfsr[92]^lfsr[113]^lfsr[115]^lfsr[117]^lfsr[119];
  assign  o_lfsr[211] = lfsr[40]^lfsr[44]^lfsr[85]^lfsr[87]^lfsr[89]^lfsr[91]^lfsr[112]^lfsr[114]^lfsr[116]^lfsr[118];
  assign  o_lfsr[212] = lfsr[39]^lfsr[43]^lfsr[84]^lfsr[86]^lfsr[88]^lfsr[90]^lfsr[111]^lfsr[113]^lfsr[115]^lfsr[117];
  assign  o_lfsr[213] = lfsr[38]^lfsr[42]^lfsr[83]^lfsr[85]^lfsr[87]^lfsr[89]^lfsr[110]^lfsr[112]^lfsr[114]^lfsr[116];
  assign  o_lfsr[214] = lfsr[37]^lfsr[41]^lfsr[82]^lfsr[84]^lfsr[86]^lfsr[88]^lfsr[109]^lfsr[111]^lfsr[113]^lfsr[115];
  assign  o_lfsr[215] = lfsr[36]^lfsr[40]^lfsr[81]^lfsr[83]^lfsr[85]^lfsr[87]^lfsr[108]^lfsr[110]^lfsr[112]^lfsr[114];
  assign  o_lfsr[216] = lfsr[35]^lfsr[39]^lfsr[80]^lfsr[82]^lfsr[84]^lfsr[86]^lfsr[107]^lfsr[109]^lfsr[111]^lfsr[113];
  assign  o_lfsr[217] = lfsr[34]^lfsr[38]^lfsr[79]^lfsr[81]^lfsr[83]^lfsr[85]^lfsr[106]^lfsr[108]^lfsr[110]^lfsr[112];
  assign  o_lfsr[218] = lfsr[33]^lfsr[37]^lfsr[78]^lfsr[80]^lfsr[82]^lfsr[84]^lfsr[105]^lfsr[107]^lfsr[109]^lfsr[111];
  assign  o_lfsr[219] = lfsr[32]^lfsr[36]^lfsr[77]^lfsr[79]^lfsr[81]^lfsr[83]^lfsr[104]^lfsr[106]^lfsr[108]^lfsr[110];
  assign  o_lfsr[220] = lfsr[31]^lfsr[35]^lfsr[76]^lfsr[78]^lfsr[80]^lfsr[82]^lfsr[103]^lfsr[105]^lfsr[107]^lfsr[109];
  assign  o_lfsr[221] = lfsr[30]^lfsr[34]^lfsr[75]^lfsr[77]^lfsr[79]^lfsr[81]^lfsr[102]^lfsr[104]^lfsr[106]^lfsr[108];
  assign  o_lfsr[222] = lfsr[29]^lfsr[33]^lfsr[74]^lfsr[76]^lfsr[78]^lfsr[80]^lfsr[101]^lfsr[103]^lfsr[105]^lfsr[107];
  assign  o_lfsr[223] = lfsr[28]^lfsr[32]^lfsr[73]^lfsr[75]^lfsr[77]^lfsr[79]^lfsr[100]^lfsr[102]^lfsr[104]^lfsr[106];
  assign  o_lfsr[224] = lfsr[27]^lfsr[31]^lfsr[72]^lfsr[74]^lfsr[76]^lfsr[78]^lfsr[99]^lfsr[101]^lfsr[103]^lfsr[105];
  assign  o_lfsr[225] = lfsr[26]^lfsr[30]^lfsr[71]^lfsr[73]^lfsr[75]^lfsr[77]^lfsr[98]^lfsr[100]^lfsr[102]^lfsr[104];
  assign  o_lfsr[226] = lfsr[25]^lfsr[29]^lfsr[70]^lfsr[72]^lfsr[74]^lfsr[76]^lfsr[97]^lfsr[99]^lfsr[101]^lfsr[103];
  assign  o_lfsr[227] = lfsr[24]^lfsr[28]^lfsr[69]^lfsr[71]^lfsr[73]^lfsr[75]^lfsr[96]^lfsr[98]^lfsr[100]^lfsr[102];
  assign  o_lfsr[228] = lfsr[23]^lfsr[27]^lfsr[68]^lfsr[70]^lfsr[72]^lfsr[74]^lfsr[95]^lfsr[97]^lfsr[99]^lfsr[101];
  assign  o_lfsr[229] = lfsr[22]^lfsr[26]^lfsr[67]^lfsr[69]^lfsr[71]^lfsr[73]^lfsr[94]^lfsr[96]^lfsr[98]^lfsr[100];
  assign  o_lfsr[230] = lfsr[21]^lfsr[25]^lfsr[66]^lfsr[68]^lfsr[70]^lfsr[72]^lfsr[93]^lfsr[95]^lfsr[97]^lfsr[99];
  assign  o_lfsr[231] = lfsr[20]^lfsr[24]^lfsr[65]^lfsr[67]^lfsr[69]^lfsr[71]^lfsr[92]^lfsr[94]^lfsr[96]^lfsr[98];
  assign  o_lfsr[232] = lfsr[19]^lfsr[23]^lfsr[64]^lfsr[66]^lfsr[68]^lfsr[70]^lfsr[91]^lfsr[93]^lfsr[95]^lfsr[97];
  assign  o_lfsr[233] = lfsr[18]^lfsr[22]^lfsr[63]^lfsr[65]^lfsr[67]^lfsr[69]^lfsr[90]^lfsr[92]^lfsr[94]^lfsr[96];
  assign  o_lfsr[234] = lfsr[17]^lfsr[21]^lfsr[62]^lfsr[64]^lfsr[66]^lfsr[68]^lfsr[89]^lfsr[91]^lfsr[93]^lfsr[95];
  assign  o_lfsr[235] = lfsr[16]^lfsr[20]^lfsr[61]^lfsr[63]^lfsr[65]^lfsr[67]^lfsr[88]^lfsr[90]^lfsr[92]^lfsr[94];
  assign  o_lfsr[236] = lfsr[15]^lfsr[19]^lfsr[60]^lfsr[62]^lfsr[64]^lfsr[66]^lfsr[87]^lfsr[89]^lfsr[91]^lfsr[93];
  assign  o_lfsr[237] = lfsr[14]^lfsr[18]^lfsr[59]^lfsr[61]^lfsr[63]^lfsr[65]^lfsr[86]^lfsr[88]^lfsr[90]^lfsr[92];
  assign  o_lfsr[238] = lfsr[13]^lfsr[17]^lfsr[58]^lfsr[60]^lfsr[62]^lfsr[64]^lfsr[85]^lfsr[87]^lfsr[89]^lfsr[91];
  assign  o_lfsr[239] = lfsr[12]^lfsr[16]^lfsr[57]^lfsr[59]^lfsr[61]^lfsr[63]^lfsr[84]^lfsr[86]^lfsr[88]^lfsr[90];
  assign  o_lfsr[240] = lfsr[11]^lfsr[15]^lfsr[56]^lfsr[58]^lfsr[60]^lfsr[62]^lfsr[83]^lfsr[85]^lfsr[87]^lfsr[89];
  assign  o_lfsr[241] = lfsr[10]^lfsr[14]^lfsr[55]^lfsr[57]^lfsr[59]^lfsr[61]^lfsr[82]^lfsr[84]^lfsr[86]^lfsr[88];
  assign  o_lfsr[242] = lfsr[ 9]^lfsr[13]^lfsr[54]^lfsr[56]^lfsr[58]^lfsr[60]^lfsr[81]^lfsr[83]^lfsr[85]^lfsr[87];
  assign  o_lfsr[243] = lfsr[ 8]^lfsr[12]^lfsr[53]^lfsr[55]^lfsr[57]^lfsr[59]^lfsr[80]^lfsr[82]^lfsr[84]^lfsr[86];
  assign  o_lfsr[244] = lfsr[ 7]^lfsr[11]^lfsr[52]^lfsr[54]^lfsr[56]^lfsr[58]^lfsr[79]^lfsr[81]^lfsr[83]^lfsr[85];
  assign  o_lfsr[245] = lfsr[ 6]^lfsr[10]^lfsr[51]^lfsr[53]^lfsr[55]^lfsr[57]^lfsr[78]^lfsr[80]^lfsr[82]^lfsr[84];
  assign  o_lfsr[246] = lfsr[ 5]^lfsr[ 9]^lfsr[50]^lfsr[52]^lfsr[54]^lfsr[56]^lfsr[77]^lfsr[79]^lfsr[81]^lfsr[83];
  assign  o_lfsr[247] = lfsr[ 4]^lfsr[ 8]^lfsr[49]^lfsr[51]^lfsr[53]^lfsr[55]^lfsr[76]^lfsr[78]^lfsr[80]^lfsr[82];
  assign  o_lfsr[248] = lfsr[ 3]^lfsr[ 7]^lfsr[48]^lfsr[50]^lfsr[52]^lfsr[54]^lfsr[75]^lfsr[77]^lfsr[79]^lfsr[81];
  assign  o_lfsr[249] = lfsr[ 2]^lfsr[ 6]^lfsr[47]^lfsr[49]^lfsr[51]^lfsr[53]^lfsr[74]^lfsr[76]^lfsr[78]^lfsr[80];
  assign  o_lfsr[250] = lfsr[ 1]^lfsr[ 5]^lfsr[46]^lfsr[48]^lfsr[50]^lfsr[52]^lfsr[73]^lfsr[75]^lfsr[77]^lfsr[79];
  assign  o_lfsr[251] = lfsr[ 0]^lfsr[ 4]^lfsr[45]^lfsr[47]^lfsr[49]^lfsr[51]^lfsr[72]^lfsr[74]^lfsr[76]^lfsr[78];
  assign  o_lfsr[252] = lfsr[ 3]^lfsr[44]^lfsr[46]^lfsr[48]^lfsr[50]^lfsr[71]^lfsr[73]^lfsr[75]^lfsr[77]^lfsr[98]^lfsr[100]^lfsr[125]^lfsr[127];
  assign  o_lfsr[253] = lfsr[ 2]^lfsr[43]^lfsr[45]^lfsr[47]^lfsr[49]^lfsr[70]^lfsr[72]^lfsr[74]^lfsr[76]^lfsr[97]^lfsr[99]^lfsr[124]^lfsr[126];
  assign  o_lfsr[254] = lfsr[ 1]^lfsr[42]^lfsr[44]^lfsr[46]^lfsr[48]^lfsr[69]^lfsr[71]^lfsr[73]^lfsr[75]^lfsr[96]^lfsr[98]^lfsr[123]^lfsr[125];
  assign  o_lfsr[255] = lfsr[ 0]^lfsr[41]^lfsr[43]^lfsr[45]^lfsr[47]^lfsr[68]^lfsr[70]^lfsr[72]^lfsr[74]^lfsr[95]^lfsr[97]^lfsr[122]^lfsr[124];
  assign  o_lfsr[256] = lfsr[40]^lfsr[42]^lfsr[44]^lfsr[46]^lfsr[67]^lfsr[69]^lfsr[71]^lfsr[73]^lfsr[94]^lfsr[96]^lfsr[98]^lfsr[100]^lfsr[121]^lfsr[123]^lfsr[125]^lfsr[127];
  assign  o_lfsr[257] = lfsr[39]^lfsr[41]^lfsr[43]^lfsr[45]^lfsr[66]^lfsr[68]^lfsr[70]^lfsr[72]^lfsr[93]^lfsr[95]^lfsr[97]^lfsr[99]^lfsr[120]^lfsr[122]^lfsr[124]^lfsr[126];
  assign  o_lfsr[258] = lfsr[38]^lfsr[40]^lfsr[42]^lfsr[44]^lfsr[65]^lfsr[67]^lfsr[69]^lfsr[71]^lfsr[92]^lfsr[94]^lfsr[96]^lfsr[98]^lfsr[119]^lfsr[121]^lfsr[123]^lfsr[125];
  assign  o_lfsr[259] = lfsr[37]^lfsr[39]^lfsr[41]^lfsr[43]^lfsr[64]^lfsr[66]^lfsr[68]^lfsr[70]^lfsr[91]^lfsr[93]^lfsr[95]^lfsr[97]^lfsr[118]^lfsr[120]^lfsr[122]^lfsr[124];
  assign  o_lfsr[260] = lfsr[36]^lfsr[38]^lfsr[40]^lfsr[42]^lfsr[63]^lfsr[65]^lfsr[67]^lfsr[69]^lfsr[90]^lfsr[92]^lfsr[94]^lfsr[96]^lfsr[117]^lfsr[119]^lfsr[121]^lfsr[123];
  assign  o_lfsr[261] = lfsr[35]^lfsr[37]^lfsr[39]^lfsr[41]^lfsr[62]^lfsr[64]^lfsr[66]^lfsr[68]^lfsr[89]^lfsr[91]^lfsr[93]^lfsr[95]^lfsr[116]^lfsr[118]^lfsr[120]^lfsr[122];
  assign  o_lfsr[262] = lfsr[34]^lfsr[36]^lfsr[38]^lfsr[40]^lfsr[61]^lfsr[63]^lfsr[65]^lfsr[67]^lfsr[88]^lfsr[90]^lfsr[92]^lfsr[94]^lfsr[115]^lfsr[117]^lfsr[119]^lfsr[121];
  assign  o_lfsr[263] = lfsr[33]^lfsr[35]^lfsr[37]^lfsr[39]^lfsr[60]^lfsr[62]^lfsr[64]^lfsr[66]^lfsr[87]^lfsr[89]^lfsr[91]^lfsr[93]^lfsr[114]^lfsr[116]^lfsr[118]^lfsr[120];
  assign  o_lfsr[264] = lfsr[32]^lfsr[34]^lfsr[36]^lfsr[38]^lfsr[59]^lfsr[61]^lfsr[63]^lfsr[65]^lfsr[86]^lfsr[88]^lfsr[90]^lfsr[92]^lfsr[113]^lfsr[115]^lfsr[117]^lfsr[119];
  assign  o_lfsr[265] = lfsr[31]^lfsr[33]^lfsr[35]^lfsr[37]^lfsr[58]^lfsr[60]^lfsr[62]^lfsr[64]^lfsr[85]^lfsr[87]^lfsr[89]^lfsr[91]^lfsr[112]^lfsr[114]^lfsr[116]^lfsr[118];
  assign  o_lfsr[266] = lfsr[30]^lfsr[32]^lfsr[34]^lfsr[36]^lfsr[57]^lfsr[59]^lfsr[61]^lfsr[63]^lfsr[84]^lfsr[86]^lfsr[88]^lfsr[90]^lfsr[111]^lfsr[113]^lfsr[115]^lfsr[117];
  assign  o_lfsr[267] = lfsr[29]^lfsr[31]^lfsr[33]^lfsr[35]^lfsr[56]^lfsr[58]^lfsr[60]^lfsr[62]^lfsr[83]^lfsr[85]^lfsr[87]^lfsr[89]^lfsr[110]^lfsr[112]^lfsr[114]^lfsr[116];
  assign  o_lfsr[268] = lfsr[28]^lfsr[30]^lfsr[32]^lfsr[34]^lfsr[55]^lfsr[57]^lfsr[59]^lfsr[61]^lfsr[82]^lfsr[84]^lfsr[86]^lfsr[88]^lfsr[109]^lfsr[111]^lfsr[113]^lfsr[115];
  assign  o_lfsr[269] = lfsr[27]^lfsr[29]^lfsr[31]^lfsr[33]^lfsr[54]^lfsr[56]^lfsr[58]^lfsr[60]^lfsr[81]^lfsr[83]^lfsr[85]^lfsr[87]^lfsr[108]^lfsr[110]^lfsr[112]^lfsr[114];
  assign  o_lfsr[270] = lfsr[26]^lfsr[28]^lfsr[30]^lfsr[32]^lfsr[53]^lfsr[55]^lfsr[57]^lfsr[59]^lfsr[80]^lfsr[82]^lfsr[84]^lfsr[86]^lfsr[107]^lfsr[109]^lfsr[111]^lfsr[113];
  assign  o_lfsr[271] = lfsr[25]^lfsr[27]^lfsr[29]^lfsr[31]^lfsr[52]^lfsr[54]^lfsr[56]^lfsr[58]^lfsr[79]^lfsr[81]^lfsr[83]^lfsr[85]^lfsr[106]^lfsr[108]^lfsr[110]^lfsr[112];
  assign  o_lfsr[272] = lfsr[24]^lfsr[26]^lfsr[28]^lfsr[30]^lfsr[51]^lfsr[53]^lfsr[55]^lfsr[57]^lfsr[78]^lfsr[80]^lfsr[82]^lfsr[84]^lfsr[105]^lfsr[107]^lfsr[109]^lfsr[111];
  assign  o_lfsr[273] = lfsr[23]^lfsr[25]^lfsr[27]^lfsr[29]^lfsr[50]^lfsr[52]^lfsr[54]^lfsr[56]^lfsr[77]^lfsr[79]^lfsr[81]^lfsr[83]^lfsr[104]^lfsr[106]^lfsr[108]^lfsr[110];
  assign  o_lfsr[274] = lfsr[22]^lfsr[24]^lfsr[26]^lfsr[28]^lfsr[49]^lfsr[51]^lfsr[53]^lfsr[55]^lfsr[76]^lfsr[78]^lfsr[80]^lfsr[82]^lfsr[103]^lfsr[105]^lfsr[107]^lfsr[109];
  assign  o_lfsr[275] = lfsr[21]^lfsr[23]^lfsr[25]^lfsr[27]^lfsr[48]^lfsr[50]^lfsr[52]^lfsr[54]^lfsr[75]^lfsr[77]^lfsr[79]^lfsr[81]^lfsr[102]^lfsr[104]^lfsr[106]^lfsr[108];
  assign  o_lfsr[276] = lfsr[20]^lfsr[22]^lfsr[24]^lfsr[26]^lfsr[47]^lfsr[49]^lfsr[51]^lfsr[53]^lfsr[74]^lfsr[76]^lfsr[78]^lfsr[80]^lfsr[101]^lfsr[103]^lfsr[105]^lfsr[107];
  assign  o_lfsr[277] = lfsr[19]^lfsr[21]^lfsr[23]^lfsr[25]^lfsr[46]^lfsr[48]^lfsr[50]^lfsr[52]^lfsr[73]^lfsr[75]^lfsr[77]^lfsr[79]^lfsr[100]^lfsr[102]^lfsr[104]^lfsr[106];
  assign  o_lfsr[278] = lfsr[18]^lfsr[20]^lfsr[22]^lfsr[24]^lfsr[45]^lfsr[47]^lfsr[49]^lfsr[51]^lfsr[72]^lfsr[74]^lfsr[76]^lfsr[78]^lfsr[99]^lfsr[101]^lfsr[103]^lfsr[105];
  assign  o_lfsr[279] = lfsr[17]^lfsr[19]^lfsr[21]^lfsr[23]^lfsr[44]^lfsr[46]^lfsr[48]^lfsr[50]^lfsr[71]^lfsr[73]^lfsr[75]^lfsr[77]^lfsr[98]^lfsr[100]^lfsr[102]^lfsr[104];
  assign  o_lfsr[280] = lfsr[16]^lfsr[18]^lfsr[20]^lfsr[22]^lfsr[43]^lfsr[45]^lfsr[47]^lfsr[49]^lfsr[70]^lfsr[72]^lfsr[74]^lfsr[76]^lfsr[97]^lfsr[99]^lfsr[101]^lfsr[103];
  assign  o_lfsr[281] = lfsr[15]^lfsr[17]^lfsr[19]^lfsr[21]^lfsr[42]^lfsr[44]^lfsr[46]^lfsr[48]^lfsr[69]^lfsr[71]^lfsr[73]^lfsr[75]^lfsr[96]^lfsr[98]^lfsr[100]^lfsr[102];
  assign  o_lfsr[282] = lfsr[14]^lfsr[16]^lfsr[18]^lfsr[20]^lfsr[41]^lfsr[43]^lfsr[45]^lfsr[47]^lfsr[68]^lfsr[70]^lfsr[72]^lfsr[74]^lfsr[95]^lfsr[97]^lfsr[99]^lfsr[101];
  assign  o_lfsr[283] = lfsr[13]^lfsr[15]^lfsr[17]^lfsr[19]^lfsr[40]^lfsr[42]^lfsr[44]^lfsr[46]^lfsr[67]^lfsr[69]^lfsr[71]^lfsr[73]^lfsr[94]^lfsr[96]^lfsr[98]^lfsr[100];
  assign  o_lfsr[284] = lfsr[12]^lfsr[14]^lfsr[16]^lfsr[18]^lfsr[39]^lfsr[41]^lfsr[43]^lfsr[45]^lfsr[66]^lfsr[68]^lfsr[70]^lfsr[72]^lfsr[93]^lfsr[95]^lfsr[97]^lfsr[99];
  assign  o_lfsr[285] = lfsr[11]^lfsr[13]^lfsr[15]^lfsr[17]^lfsr[38]^lfsr[40]^lfsr[42]^lfsr[44]^lfsr[65]^lfsr[67]^lfsr[69]^lfsr[71]^lfsr[92]^lfsr[94]^lfsr[96]^lfsr[98];
  assign  o_lfsr[286] = lfsr[10]^lfsr[12]^lfsr[14]^lfsr[16]^lfsr[37]^lfsr[39]^lfsr[41]^lfsr[43]^lfsr[64]^lfsr[66]^lfsr[68]^lfsr[70]^lfsr[91]^lfsr[93]^lfsr[95]^lfsr[97];
  assign  o_lfsr[287] = lfsr[ 9]^lfsr[11]^lfsr[13]^lfsr[15]^lfsr[36]^lfsr[38]^lfsr[40]^lfsr[42]^lfsr[63]^lfsr[65]^lfsr[67]^lfsr[69]^lfsr[90]^lfsr[92]^lfsr[94]^lfsr[96];
  assign  o_lfsr[288] = lfsr[ 8]^lfsr[10]^lfsr[12]^lfsr[14]^lfsr[35]^lfsr[37]^lfsr[39]^lfsr[41]^lfsr[62]^lfsr[64]^lfsr[66]^lfsr[68]^lfsr[89]^lfsr[91]^lfsr[93]^lfsr[95];
  assign  o_lfsr[289] = lfsr[ 7]^lfsr[ 9]^lfsr[11]^lfsr[13]^lfsr[34]^lfsr[36]^lfsr[38]^lfsr[40]^lfsr[61]^lfsr[63]^lfsr[65]^lfsr[67]^lfsr[88]^lfsr[90]^lfsr[92]^lfsr[94];
  assign  o_lfsr[290] = lfsr[ 6]^lfsr[ 8]^lfsr[10]^lfsr[12]^lfsr[33]^lfsr[35]^lfsr[37]^lfsr[39]^lfsr[60]^lfsr[62]^lfsr[64]^lfsr[66]^lfsr[87]^lfsr[89]^lfsr[91]^lfsr[93];
  assign  o_lfsr[291] = lfsr[ 5]^lfsr[ 7]^lfsr[ 9]^lfsr[11]^lfsr[32]^lfsr[34]^lfsr[36]^lfsr[38]^lfsr[59]^lfsr[61]^lfsr[63]^lfsr[65]^lfsr[86]^lfsr[88]^lfsr[90]^lfsr[92];
  assign  o_lfsr[292] = lfsr[ 4]^lfsr[ 6]^lfsr[ 8]^lfsr[10]^lfsr[31]^lfsr[33]^lfsr[35]^lfsr[37]^lfsr[58]^lfsr[60]^lfsr[62]^lfsr[64]^lfsr[85]^lfsr[87]^lfsr[89]^lfsr[91];
  assign  o_lfsr[293] = lfsr[ 3]^lfsr[ 5]^lfsr[ 7]^lfsr[ 9]^lfsr[30]^lfsr[32]^lfsr[34]^lfsr[36]^lfsr[57]^lfsr[59]^lfsr[61]^lfsr[63]^lfsr[84]^lfsr[86]^lfsr[88]^lfsr[90];
  assign  o_lfsr[294] = lfsr[ 2]^lfsr[ 4]^lfsr[ 6]^lfsr[ 8]^lfsr[29]^lfsr[31]^lfsr[33]^lfsr[35]^lfsr[56]^lfsr[58]^lfsr[60]^lfsr[62]^lfsr[83]^lfsr[85]^lfsr[87]^lfsr[89];
  assign  o_lfsr[295] = lfsr[ 1]^lfsr[ 3]^lfsr[ 5]^lfsr[ 7]^lfsr[28]^lfsr[30]^lfsr[32]^lfsr[34]^lfsr[55]^lfsr[57]^lfsr[59]^lfsr[61]^lfsr[82]^lfsr[84]^lfsr[86]^lfsr[88];
  assign  o_lfsr[296] = lfsr[ 0]^lfsr[ 2]^lfsr[ 4]^lfsr[ 6]^lfsr[27]^lfsr[29]^lfsr[31]^lfsr[33]^lfsr[54]^lfsr[56]^lfsr[58]^lfsr[60]^lfsr[81]^lfsr[83]^lfsr[85]^lfsr[87];
  assign  o_lfsr[297] = lfsr[ 1]^lfsr[ 3]^lfsr[ 5]^lfsr[26]^lfsr[28]^lfsr[30]^lfsr[32]^lfsr[53]^lfsr[55]^lfsr[57]^lfsr[59]^lfsr[80]^lfsr[82]^lfsr[84]^lfsr[86]^lfsr[98]^lfsr[100]^lfsr[125]^lfsr[127];
  assign  o_lfsr[298] = lfsr[ 0]^lfsr[ 2]^lfsr[ 4]^lfsr[25]^lfsr[27]^lfsr[29]^lfsr[31]^lfsr[52]^lfsr[54]^lfsr[56]^lfsr[58]^lfsr[79]^lfsr[81]^lfsr[83]^lfsr[85]^lfsr[97]^lfsr[99]^lfsr[124]^lfsr[126];
  assign  o_lfsr[299] = lfsr[ 1]^lfsr[ 3]^lfsr[24]^lfsr[26]^lfsr[28]^lfsr[30]^lfsr[51]^lfsr[53]^lfsr[55]^lfsr[57]^lfsr[78]^lfsr[80]^lfsr[82]^lfsr[84]^lfsr[96]^lfsr[100]^lfsr[123]^lfsr[127];
  assign  o_lfsr[300] = lfsr[ 0]^lfsr[ 2]^lfsr[23]^lfsr[25]^lfsr[27]^lfsr[29]^lfsr[50]^lfsr[52]^lfsr[54]^lfsr[56]^lfsr[77]^lfsr[79]^lfsr[81]^lfsr[83]^lfsr[95]^lfsr[99]^lfsr[122]^lfsr[126];
  assign  o_lfsr[301] = lfsr[ 1]^lfsr[22]^lfsr[24]^lfsr[26]^lfsr[28]^lfsr[49]^lfsr[51]^lfsr[53]^lfsr[55]^lfsr[76]^lfsr[78]^lfsr[80]^lfsr[82]^lfsr[94]^lfsr[100]^lfsr[121]^lfsr[127];
  assign  o_lfsr[302] = lfsr[ 0]^lfsr[21]^lfsr[23]^lfsr[25]^lfsr[27]^lfsr[48]^lfsr[50]^lfsr[52]^lfsr[54]^lfsr[75]^lfsr[77]^lfsr[79]^lfsr[81]^lfsr[93]^lfsr[99]^lfsr[120]^lfsr[126];
  assign  o_lfsr[303] = lfsr[20]^lfsr[22]^lfsr[24]^lfsr[26]^lfsr[47]^lfsr[49]^lfsr[51]^lfsr[53]^lfsr[74]^lfsr[76]^lfsr[78]^lfsr[80]^lfsr[92]^lfsr[100]^lfsr[119]^lfsr[127];
  assign  o_lfsr[304] = lfsr[19]^lfsr[21]^lfsr[23]^lfsr[25]^lfsr[46]^lfsr[48]^lfsr[50]^lfsr[52]^lfsr[73]^lfsr[75]^lfsr[77]^lfsr[79]^lfsr[91]^lfsr[99]^lfsr[118]^lfsr[126];
  assign  o_lfsr[305] = lfsr[18]^lfsr[20]^lfsr[22]^lfsr[24]^lfsr[45]^lfsr[47]^lfsr[49]^lfsr[51]^lfsr[72]^lfsr[74]^lfsr[76]^lfsr[78]^lfsr[90]^lfsr[98]^lfsr[117]^lfsr[125];
  assign  o_lfsr[306] = lfsr[17]^lfsr[19]^lfsr[21]^lfsr[23]^lfsr[44]^lfsr[46]^lfsr[48]^lfsr[50]^lfsr[71]^lfsr[73]^lfsr[75]^lfsr[77]^lfsr[89]^lfsr[97]^lfsr[116]^lfsr[124];
  assign  o_lfsr[307] = lfsr[16]^lfsr[18]^lfsr[20]^lfsr[22]^lfsr[43]^lfsr[45]^lfsr[47]^lfsr[49]^lfsr[70]^lfsr[72]^lfsr[74]^lfsr[76]^lfsr[88]^lfsr[96]^lfsr[115]^lfsr[123];
  assign  o_lfsr[308] = lfsr[15]^lfsr[17]^lfsr[19]^lfsr[21]^lfsr[42]^lfsr[44]^lfsr[46]^lfsr[48]^lfsr[69]^lfsr[71]^lfsr[73]^lfsr[75]^lfsr[87]^lfsr[95]^lfsr[114]^lfsr[122];
  assign  o_lfsr[309] = lfsr[14]^lfsr[16]^lfsr[18]^lfsr[20]^lfsr[41]^lfsr[43]^lfsr[45]^lfsr[47]^lfsr[68]^lfsr[70]^lfsr[72]^lfsr[74]^lfsr[86]^lfsr[94]^lfsr[113]^lfsr[121];
  assign  o_lfsr[310] = lfsr[13]^lfsr[15]^lfsr[17]^lfsr[19]^lfsr[40]^lfsr[42]^lfsr[44]^lfsr[46]^lfsr[67]^lfsr[69]^lfsr[71]^lfsr[73]^lfsr[85]^lfsr[93]^lfsr[112]^lfsr[120];
  assign  o_lfsr[311] = lfsr[12]^lfsr[14]^lfsr[16]^lfsr[18]^lfsr[39]^lfsr[41]^lfsr[43]^lfsr[45]^lfsr[66]^lfsr[68]^lfsr[70]^lfsr[72]^lfsr[84]^lfsr[92]^lfsr[111]^lfsr[119];
  assign  o_lfsr[312] = lfsr[11]^lfsr[13]^lfsr[15]^lfsr[17]^lfsr[38]^lfsr[40]^lfsr[42]^lfsr[44]^lfsr[65]^lfsr[67]^lfsr[69]^lfsr[71]^lfsr[83]^lfsr[91]^lfsr[110]^lfsr[118];
  assign  o_lfsr[313] = lfsr[10]^lfsr[12]^lfsr[14]^lfsr[16]^lfsr[37]^lfsr[39]^lfsr[41]^lfsr[43]^lfsr[64]^lfsr[66]^lfsr[68]^lfsr[70]^lfsr[82]^lfsr[90]^lfsr[109]^lfsr[117];
  assign  o_lfsr[314] = lfsr[ 9]^lfsr[11]^lfsr[13]^lfsr[15]^lfsr[36]^lfsr[38]^lfsr[40]^lfsr[42]^lfsr[63]^lfsr[65]^lfsr[67]^lfsr[69]^lfsr[81]^lfsr[89]^lfsr[108]^lfsr[116];
  assign  o_lfsr[315] = lfsr[ 8]^lfsr[10]^lfsr[12]^lfsr[14]^lfsr[35]^lfsr[37]^lfsr[39]^lfsr[41]^lfsr[62]^lfsr[64]^lfsr[66]^lfsr[68]^lfsr[80]^lfsr[88]^lfsr[107]^lfsr[115];
  assign  o_lfsr[316] = lfsr[ 7]^lfsr[ 9]^lfsr[11]^lfsr[13]^lfsr[34]^lfsr[36]^lfsr[38]^lfsr[40]^lfsr[61]^lfsr[63]^lfsr[65]^lfsr[67]^lfsr[79]^lfsr[87]^lfsr[106]^lfsr[114];
  assign  o_lfsr[317] = lfsr[ 6]^lfsr[ 8]^lfsr[10]^lfsr[12]^lfsr[33]^lfsr[35]^lfsr[37]^lfsr[39]^lfsr[60]^lfsr[62]^lfsr[64]^lfsr[66]^lfsr[78]^lfsr[86]^lfsr[105]^lfsr[113];
  assign  o_lfsr[318] = lfsr[ 5]^lfsr[ 7]^lfsr[ 9]^lfsr[11]^lfsr[32]^lfsr[34]^lfsr[36]^lfsr[38]^lfsr[59]^lfsr[61]^lfsr[63]^lfsr[65]^lfsr[77]^lfsr[85]^lfsr[104]^lfsr[112];
  assign  o_lfsr[319] = lfsr[ 4]^lfsr[ 6]^lfsr[ 8]^lfsr[10]^lfsr[31]^lfsr[33]^lfsr[35]^lfsr[37]^lfsr[58]^lfsr[60]^lfsr[62]^lfsr[64]^lfsr[76]^lfsr[84]^lfsr[103]^lfsr[111];
  assign  o_lfsr[320] = lfsr[ 3]^lfsr[ 5]^lfsr[ 7]^lfsr[ 9]^lfsr[30]^lfsr[32]^lfsr[34]^lfsr[36]^lfsr[57]^lfsr[59]^lfsr[61]^lfsr[63]^lfsr[75]^lfsr[83]^lfsr[102]^lfsr[110];
  assign  o_lfsr[321] = lfsr[ 2]^lfsr[ 4]^lfsr[ 6]^lfsr[ 8]^lfsr[29]^lfsr[31]^lfsr[33]^lfsr[35]^lfsr[56]^lfsr[58]^lfsr[60]^lfsr[62]^lfsr[74]^lfsr[82]^lfsr[101]^lfsr[109];
  assign  o_lfsr[322] = lfsr[ 1]^lfsr[ 3]^lfsr[ 5]^lfsr[ 7]^lfsr[28]^lfsr[30]^lfsr[32]^lfsr[34]^lfsr[55]^lfsr[57]^lfsr[59]^lfsr[61]^lfsr[73]^lfsr[81]^lfsr[100]^lfsr[108];
  assign  o_lfsr[323] = lfsr[ 0]^lfsr[ 2]^lfsr[ 4]^lfsr[ 6]^lfsr[27]^lfsr[29]^lfsr[31]^lfsr[33]^lfsr[54]^lfsr[56]^lfsr[58]^lfsr[60]^lfsr[72]^lfsr[80]^lfsr[99]^lfsr[107];
  assign  o_lfsr[324] = lfsr[ 1]^lfsr[ 3]^lfsr[ 5]^lfsr[26]^lfsr[28]^lfsr[30]^lfsr[32]^lfsr[53]^lfsr[55]^lfsr[57]^lfsr[59]^lfsr[71]^lfsr[79]^lfsr[100]^lfsr[106]^lfsr[125]^lfsr[127];
  assign  o_lfsr[325] = lfsr[ 0]^lfsr[ 2]^lfsr[ 4]^lfsr[25]^lfsr[27]^lfsr[29]^lfsr[31]^lfsr[52]^lfsr[54]^lfsr[56]^lfsr[58]^lfsr[70]^lfsr[78]^lfsr[99]^lfsr[105]^lfsr[124]^lfsr[126];
  assign  o_lfsr[326] = lfsr[ 1]^lfsr[ 3]^lfsr[24]^lfsr[26]^lfsr[28]^lfsr[30]^lfsr[51]^lfsr[53]^lfsr[55]^lfsr[57]^lfsr[69]^lfsr[77]^lfsr[100]^lfsr[104]^lfsr[123]^lfsr[127];
  assign  o_lfsr[327] = lfsr[ 0]^lfsr[ 2]^lfsr[23]^lfsr[25]^lfsr[27]^lfsr[29]^lfsr[50]^lfsr[52]^lfsr[54]^lfsr[56]^lfsr[68]^lfsr[76]^lfsr[99]^lfsr[103]^lfsr[122]^lfsr[126];
  assign  o_lfsr[328] = lfsr[ 1]^lfsr[22]^lfsr[24]^lfsr[26]^lfsr[28]^lfsr[49]^lfsr[51]^lfsr[53]^lfsr[55]^lfsr[67]^lfsr[75]^lfsr[100]^lfsr[102]^lfsr[121]^lfsr[127];
  assign  o_lfsr[329] = lfsr[ 0]^lfsr[21]^lfsr[23]^lfsr[25]^lfsr[27]^lfsr[48]^lfsr[50]^lfsr[52]^lfsr[54]^lfsr[66]^lfsr[74]^lfsr[99]^lfsr[101]^lfsr[120]^lfsr[126];
  assign  o_lfsr[330] = lfsr[20]^lfsr[22]^lfsr[24]^lfsr[26]^lfsr[47]^lfsr[49]^lfsr[51]^lfsr[53]^lfsr[65]^lfsr[73]^lfsr[119]^lfsr[127];
  assign  o_lfsr[331] = lfsr[19]^lfsr[21]^lfsr[23]^lfsr[25]^lfsr[46]^lfsr[48]^lfsr[50]^lfsr[52]^lfsr[64]^lfsr[72]^lfsr[118]^lfsr[126];
  assign  o_lfsr[332] = lfsr[18]^lfsr[20]^lfsr[22]^lfsr[24]^lfsr[45]^lfsr[47]^lfsr[49]^lfsr[51]^lfsr[63]^lfsr[71]^lfsr[117]^lfsr[125];
  assign  o_lfsr[333] = lfsr[17]^lfsr[19]^lfsr[21]^lfsr[23]^lfsr[44]^lfsr[46]^lfsr[48]^lfsr[50]^lfsr[62]^lfsr[70]^lfsr[116]^lfsr[124];
  assign  o_lfsr[334] = lfsr[16]^lfsr[18]^lfsr[20]^lfsr[22]^lfsr[43]^lfsr[45]^lfsr[47]^lfsr[49]^lfsr[61]^lfsr[69]^lfsr[115]^lfsr[123];
  assign  o_lfsr[335] = lfsr[15]^lfsr[17]^lfsr[19]^lfsr[21]^lfsr[42]^lfsr[44]^lfsr[46]^lfsr[48]^lfsr[60]^lfsr[68]^lfsr[114]^lfsr[122];
  assign  o_lfsr[336] = lfsr[14]^lfsr[16]^lfsr[18]^lfsr[20]^lfsr[41]^lfsr[43]^lfsr[45]^lfsr[47]^lfsr[59]^lfsr[67]^lfsr[113]^lfsr[121];
  assign  o_lfsr[337] = lfsr[13]^lfsr[15]^lfsr[17]^lfsr[19]^lfsr[40]^lfsr[42]^lfsr[44]^lfsr[46]^lfsr[58]^lfsr[66]^lfsr[112]^lfsr[120];
  assign  o_lfsr[338] = lfsr[12]^lfsr[14]^lfsr[16]^lfsr[18]^lfsr[39]^lfsr[41]^lfsr[43]^lfsr[45]^lfsr[57]^lfsr[65]^lfsr[111]^lfsr[119];
  assign  o_lfsr[339] = lfsr[11]^lfsr[13]^lfsr[15]^lfsr[17]^lfsr[38]^lfsr[40]^lfsr[42]^lfsr[44]^lfsr[56]^lfsr[64]^lfsr[110]^lfsr[118];
  assign  o_lfsr[340] = lfsr[10]^lfsr[12]^lfsr[14]^lfsr[16]^lfsr[37]^lfsr[39]^lfsr[41]^lfsr[43]^lfsr[55]^lfsr[63]^lfsr[109]^lfsr[117];
  assign  o_lfsr[341] = lfsr[ 9]^lfsr[11]^lfsr[13]^lfsr[15]^lfsr[36]^lfsr[38]^lfsr[40]^lfsr[42]^lfsr[54]^lfsr[62]^lfsr[108]^lfsr[116];
  assign  o_lfsr[342] = lfsr[ 8]^lfsr[10]^lfsr[12]^lfsr[14]^lfsr[35]^lfsr[37]^lfsr[39]^lfsr[41]^lfsr[53]^lfsr[61]^lfsr[107]^lfsr[115];
  assign  o_lfsr[343] = lfsr[ 7]^lfsr[ 9]^lfsr[11]^lfsr[13]^lfsr[34]^lfsr[36]^lfsr[38]^lfsr[40]^lfsr[52]^lfsr[60]^lfsr[106]^lfsr[114];
  assign  o_lfsr[344] = lfsr[ 6]^lfsr[ 8]^lfsr[10]^lfsr[12]^lfsr[33]^lfsr[35]^lfsr[37]^lfsr[39]^lfsr[51]^lfsr[59]^lfsr[105]^lfsr[113];
  assign  o_lfsr[345] = lfsr[ 5]^lfsr[ 7]^lfsr[ 9]^lfsr[11]^lfsr[32]^lfsr[34]^lfsr[36]^lfsr[38]^lfsr[50]^lfsr[58]^lfsr[104]^lfsr[112];
  assign  o_lfsr[346] = lfsr[ 4]^lfsr[ 6]^lfsr[ 8]^lfsr[10]^lfsr[31]^lfsr[33]^lfsr[35]^lfsr[37]^lfsr[49]^lfsr[57]^lfsr[103]^lfsr[111];
  assign  o_lfsr[347] = lfsr[ 3]^lfsr[ 5]^lfsr[ 7]^lfsr[ 9]^lfsr[30]^lfsr[32]^lfsr[34]^lfsr[36]^lfsr[48]^lfsr[56]^lfsr[102]^lfsr[110];
  assign  o_lfsr[348] = lfsr[ 2]^lfsr[ 4]^lfsr[ 6]^lfsr[ 8]^lfsr[29]^lfsr[31]^lfsr[33]^lfsr[35]^lfsr[47]^lfsr[55]^lfsr[101]^lfsr[109];
  assign  o_lfsr[349] = lfsr[ 1]^lfsr[ 3]^lfsr[ 5]^lfsr[ 7]^lfsr[28]^lfsr[30]^lfsr[32]^lfsr[34]^lfsr[46]^lfsr[54]^lfsr[100]^lfsr[108];
  assign  o_lfsr[350] = lfsr[ 0]^lfsr[ 2]^lfsr[ 4]^lfsr[ 6]^lfsr[27]^lfsr[29]^lfsr[31]^lfsr[33]^lfsr[45]^lfsr[53]^lfsr[99]^lfsr[107];
  assign  o_lfsr[351] = lfsr[ 1]^lfsr[ 3]^lfsr[ 5]^lfsr[26]^lfsr[28]^lfsr[30]^lfsr[32]^lfsr[44]^lfsr[52]^lfsr[100]^lfsr[106]^lfsr[125]^lfsr[127];
  assign  o_lfsr[352] = lfsr[ 0]^lfsr[ 2]^lfsr[ 4]^lfsr[25]^lfsr[27]^lfsr[29]^lfsr[31]^lfsr[43]^lfsr[51]^lfsr[99]^lfsr[105]^lfsr[124]^lfsr[126];
  assign  o_lfsr[353] = lfsr[ 1]^lfsr[ 3]^lfsr[24]^lfsr[26]^lfsr[28]^lfsr[30]^lfsr[42]^lfsr[50]^lfsr[100]^lfsr[104]^lfsr[123]^lfsr[127];
  assign  o_lfsr[354] = lfsr[ 0]^lfsr[ 2]^lfsr[23]^lfsr[25]^lfsr[27]^lfsr[29]^lfsr[41]^lfsr[49]^lfsr[99]^lfsr[103]^lfsr[122]^lfsr[126];
  assign  o_lfsr[355] = lfsr[ 1]^lfsr[22]^lfsr[24]^lfsr[26]^lfsr[28]^lfsr[40]^lfsr[48]^lfsr[100]^lfsr[102]^lfsr[121]^lfsr[127];
  assign  o_lfsr[356] = lfsr[ 0]^lfsr[21]^lfsr[23]^lfsr[25]^lfsr[27]^lfsr[39]^lfsr[47]^lfsr[99]^lfsr[101]^lfsr[120]^lfsr[126];
  assign  o_lfsr[357] = lfsr[20]^lfsr[22]^lfsr[24]^lfsr[26]^lfsr[38]^lfsr[46]^lfsr[119]^lfsr[127];
  assign  o_lfsr[358] = lfsr[19]^lfsr[21]^lfsr[23]^lfsr[25]^lfsr[37]^lfsr[45]^lfsr[118]^lfsr[126];
  assign  o_lfsr[359] = lfsr[18]^lfsr[20]^lfsr[22]^lfsr[24]^lfsr[36]^lfsr[44]^lfsr[117]^lfsr[125];
  assign  o_lfsr[360] = lfsr[17]^lfsr[19]^lfsr[21]^lfsr[23]^lfsr[35]^lfsr[43]^lfsr[116]^lfsr[124];
  assign  o_lfsr[361] = lfsr[16]^lfsr[18]^lfsr[20]^lfsr[22]^lfsr[34]^lfsr[42]^lfsr[115]^lfsr[123];
  assign  o_lfsr[362] = lfsr[15]^lfsr[17]^lfsr[19]^lfsr[21]^lfsr[33]^lfsr[41]^lfsr[114]^lfsr[122];
  assign  o_lfsr[363] = lfsr[14]^lfsr[16]^lfsr[18]^lfsr[20]^lfsr[32]^lfsr[40]^lfsr[113]^lfsr[121];
  assign  o_lfsr[364] = lfsr[13]^lfsr[15]^lfsr[17]^lfsr[19]^lfsr[31]^lfsr[39]^lfsr[112]^lfsr[120];
  assign  o_lfsr[365] = lfsr[12]^lfsr[14]^lfsr[16]^lfsr[18]^lfsr[30]^lfsr[38]^lfsr[111]^lfsr[119];
  assign  o_lfsr[366] = lfsr[11]^lfsr[13]^lfsr[15]^lfsr[17]^lfsr[29]^lfsr[37]^lfsr[110]^lfsr[118];
  assign  o_lfsr[367] = lfsr[10]^lfsr[12]^lfsr[14]^lfsr[16]^lfsr[28]^lfsr[36]^lfsr[109]^lfsr[117];
  assign  o_lfsr[368] = lfsr[ 9]^lfsr[11]^lfsr[13]^lfsr[15]^lfsr[27]^lfsr[35]^lfsr[108]^lfsr[116];
  assign  o_lfsr[369] = lfsr[ 8]^lfsr[10]^lfsr[12]^lfsr[14]^lfsr[26]^lfsr[34]^lfsr[107]^lfsr[115];
  assign  o_lfsr[370] = lfsr[ 7]^lfsr[ 9]^lfsr[11]^lfsr[13]^lfsr[25]^lfsr[33]^lfsr[106]^lfsr[114];
  assign  o_lfsr[371] = lfsr[ 6]^lfsr[ 8]^lfsr[10]^lfsr[12]^lfsr[24]^lfsr[32]^lfsr[105]^lfsr[113];
  assign  o_lfsr[372] = lfsr[ 5]^lfsr[ 7]^lfsr[ 9]^lfsr[11]^lfsr[23]^lfsr[31]^lfsr[104]^lfsr[112];
  assign  o_lfsr[373] = lfsr[ 4]^lfsr[ 6]^lfsr[ 8]^lfsr[10]^lfsr[22]^lfsr[30]^lfsr[103]^lfsr[111];
  assign  o_lfsr[374] = lfsr[ 3]^lfsr[ 5]^lfsr[ 7]^lfsr[ 9]^lfsr[21]^lfsr[29]^lfsr[102]^lfsr[110];
  assign  o_lfsr[375] = lfsr[ 2]^lfsr[ 4]^lfsr[ 6]^lfsr[ 8]^lfsr[20]^lfsr[28]^lfsr[101]^lfsr[109];
  assign  o_lfsr[376] = lfsr[ 1]^lfsr[ 3]^lfsr[ 5]^lfsr[ 7]^lfsr[19]^lfsr[27]^lfsr[100]^lfsr[108];
  assign  o_lfsr[377] = lfsr[ 0]^lfsr[ 2]^lfsr[ 4]^lfsr[ 6]^lfsr[18]^lfsr[26]^lfsr[99]^lfsr[107];
  assign  o_lfsr[378] = lfsr[ 1]^lfsr[ 3]^lfsr[ 5]^lfsr[17]^lfsr[25]^lfsr[100]^lfsr[106]^lfsr[125]^lfsr[127];
  assign  o_lfsr[379] = lfsr[ 0]^lfsr[ 2]^lfsr[ 4]^lfsr[16]^lfsr[24]^lfsr[99]^lfsr[105]^lfsr[124]^lfsr[126];
  assign  o_lfsr[380] = lfsr[ 1]^lfsr[ 3]^lfsr[15]^lfsr[23]^lfsr[100]^lfsr[104]^lfsr[123]^lfsr[127];
  assign  o_lfsr[381] = lfsr[ 0]^lfsr[ 2]^lfsr[14]^lfsr[22]^lfsr[99]^lfsr[103]^lfsr[122]^lfsr[126];
  assign  o_lfsr[382] = lfsr[ 1]^lfsr[13]^lfsr[21]^lfsr[100]^lfsr[102]^lfsr[121]^lfsr[127];
  assign  o_lfsr[383] = lfsr[ 0]^lfsr[12]^lfsr[20]^lfsr[99]^lfsr[101]^lfsr[120]^lfsr[126];
  assign  o_lfsr[384] = lfsr[11]^lfsr[19]^lfsr[119]^lfsr[127];
  assign  o_lfsr[385] = lfsr[10]^lfsr[18]^lfsr[118]^lfsr[126];
  assign  o_lfsr[386] = lfsr[ 9]^lfsr[17]^lfsr[117]^lfsr[125];
  assign  o_lfsr[387] = lfsr[ 8]^lfsr[16]^lfsr[116]^lfsr[124];
  assign  o_lfsr[388] = lfsr[ 7]^lfsr[15]^lfsr[115]^lfsr[123];
  assign  o_lfsr[389] = lfsr[ 6]^lfsr[14]^lfsr[114]^lfsr[122];
  assign  o_lfsr[390] = lfsr[ 5]^lfsr[13]^lfsr[113]^lfsr[121];
  assign  o_lfsr[391] = lfsr[ 4]^lfsr[12]^lfsr[112]^lfsr[120];
  assign  o_lfsr[392] = lfsr[ 3]^lfsr[11]^lfsr[111]^lfsr[119];
  assign  o_lfsr[393] = lfsr[ 2]^lfsr[10]^lfsr[110]^lfsr[118];
  assign  o_lfsr[394] = lfsr[ 1]^lfsr[ 9]^lfsr[109]^lfsr[117];
  assign  o_lfsr[395] = lfsr[ 0]^lfsr[ 8]^lfsr[108]^lfsr[116];
  assign  o_lfsr[396] = lfsr[ 7]^lfsr[98]^lfsr[100]^lfsr[107]^lfsr[115]^lfsr[125]^lfsr[127];
  assign  o_lfsr[397] = lfsr[ 6]^lfsr[97]^lfsr[99]^lfsr[106]^lfsr[114]^lfsr[124]^lfsr[126];
  assign  o_lfsr[398] = lfsr[ 5]^lfsr[96]^lfsr[98]^lfsr[105]^lfsr[113]^lfsr[123]^lfsr[125];
  assign  o_lfsr[399] = lfsr[ 4]^lfsr[95]^lfsr[97]^lfsr[104]^lfsr[112]^lfsr[122]^lfsr[124];
  assign  o_lfsr[400] = lfsr[ 3]^lfsr[94]^lfsr[96]^lfsr[103]^lfsr[111]^lfsr[121]^lfsr[123];
  assign  o_lfsr[401] = lfsr[ 2]^lfsr[93]^lfsr[95]^lfsr[102]^lfsr[110]^lfsr[120]^lfsr[122];
  assign  o_lfsr[402] = lfsr[ 1]^lfsr[92]^lfsr[94]^lfsr[101]^lfsr[109]^lfsr[119]^lfsr[121];
  assign  o_lfsr[403] = lfsr[ 0]^lfsr[91]^lfsr[93]^lfsr[100]^lfsr[108]^lfsr[118]^lfsr[120];
  assign  o_lfsr[404] = lfsr[90]^lfsr[92]^lfsr[98]^lfsr[99]^lfsr[100]^lfsr[107]^lfsr[117]^lfsr[119]^lfsr[125]^lfsr[127];
  assign  o_lfsr[405] = lfsr[89]^lfsr[91]^lfsr[97]^lfsr[98]^lfsr[99]^lfsr[106]^lfsr[116]^lfsr[118]^lfsr[124]^lfsr[126];
  assign  o_lfsr[406] = lfsr[88]^lfsr[90]^lfsr[96]^lfsr[97]^lfsr[98]^lfsr[105]^lfsr[115]^lfsr[117]^lfsr[123]^lfsr[125];
  assign  o_lfsr[407] = lfsr[87]^lfsr[89]^lfsr[95]^lfsr[96]^lfsr[97]^lfsr[104]^lfsr[114]^lfsr[116]^lfsr[122]^lfsr[124];
  assign  o_lfsr[408] = lfsr[86]^lfsr[88]^lfsr[94]^lfsr[95]^lfsr[96]^lfsr[103]^lfsr[113]^lfsr[115]^lfsr[121]^lfsr[123];
  assign  o_lfsr[409] = lfsr[85]^lfsr[87]^lfsr[93]^lfsr[94]^lfsr[95]^lfsr[102]^lfsr[112]^lfsr[114]^lfsr[120]^lfsr[122];
  assign  o_lfsr[410] = lfsr[84]^lfsr[86]^lfsr[92]^lfsr[93]^lfsr[94]^lfsr[101]^lfsr[111]^lfsr[113]^lfsr[119]^lfsr[121];
  assign  o_lfsr[411] = lfsr[83]^lfsr[85]^lfsr[91]^lfsr[92]^lfsr[93]^lfsr[100]^lfsr[110]^lfsr[112]^lfsr[118]^lfsr[120];
  assign  o_lfsr[412] = lfsr[82]^lfsr[84]^lfsr[90]^lfsr[91]^lfsr[92]^lfsr[99]^lfsr[109]^lfsr[111]^lfsr[117]^lfsr[119];
  assign  o_lfsr[413] = lfsr[81]^lfsr[83]^lfsr[89]^lfsr[90]^lfsr[91]^lfsr[98]^lfsr[108]^lfsr[110]^lfsr[116]^lfsr[118];
  assign  o_lfsr[414] = lfsr[80]^lfsr[82]^lfsr[88]^lfsr[89]^lfsr[90]^lfsr[97]^lfsr[107]^lfsr[109]^lfsr[115]^lfsr[117];
  assign  o_lfsr[415] = lfsr[79]^lfsr[81]^lfsr[87]^lfsr[88]^lfsr[89]^lfsr[96]^lfsr[106]^lfsr[108]^lfsr[114]^lfsr[116];
  assign  o_lfsr[416] = lfsr[78]^lfsr[80]^lfsr[86]^lfsr[87]^lfsr[88]^lfsr[95]^lfsr[105]^lfsr[107]^lfsr[113]^lfsr[115];
  assign  o_lfsr[417] = lfsr[77]^lfsr[79]^lfsr[85]^lfsr[86]^lfsr[87]^lfsr[94]^lfsr[104]^lfsr[106]^lfsr[112]^lfsr[114];
  assign  o_lfsr[418] = lfsr[76]^lfsr[78]^lfsr[84]^lfsr[85]^lfsr[86]^lfsr[93]^lfsr[103]^lfsr[105]^lfsr[111]^lfsr[113];
  assign  o_lfsr[419] = lfsr[75]^lfsr[77]^lfsr[83]^lfsr[84]^lfsr[85]^lfsr[92]^lfsr[102]^lfsr[104]^lfsr[110]^lfsr[112];
  assign  o_lfsr[420] = lfsr[74]^lfsr[76]^lfsr[82]^lfsr[83]^lfsr[84]^lfsr[91]^lfsr[101]^lfsr[103]^lfsr[109]^lfsr[111];
  assign  o_lfsr[421] = lfsr[73]^lfsr[75]^lfsr[81]^lfsr[82]^lfsr[83]^lfsr[90]^lfsr[100]^lfsr[102]^lfsr[108]^lfsr[110];
  assign  o_lfsr[422] = lfsr[72]^lfsr[74]^lfsr[80]^lfsr[81]^lfsr[82]^lfsr[89]^lfsr[99]^lfsr[101]^lfsr[107]^lfsr[109];
  assign  o_lfsr[423] = lfsr[71]^lfsr[73]^lfsr[79]^lfsr[80]^lfsr[81]^lfsr[88]^lfsr[98]^lfsr[100]^lfsr[106]^lfsr[108];
  assign  o_lfsr[424] = lfsr[70]^lfsr[72]^lfsr[78]^lfsr[79]^lfsr[80]^lfsr[87]^lfsr[97]^lfsr[99]^lfsr[105]^lfsr[107];
  assign  o_lfsr[425] = lfsr[69]^lfsr[71]^lfsr[77]^lfsr[78]^lfsr[79]^lfsr[86]^lfsr[96]^lfsr[98]^lfsr[104]^lfsr[106];
  assign  o_lfsr[426] = lfsr[68]^lfsr[70]^lfsr[76]^lfsr[77]^lfsr[78]^lfsr[85]^lfsr[95]^lfsr[97]^lfsr[103]^lfsr[105];
  assign  o_lfsr[427] = lfsr[67]^lfsr[69]^lfsr[75]^lfsr[76]^lfsr[77]^lfsr[84]^lfsr[94]^lfsr[96]^lfsr[102]^lfsr[104];
  assign  o_lfsr[428] = lfsr[66]^lfsr[68]^lfsr[74]^lfsr[75]^lfsr[76]^lfsr[83]^lfsr[93]^lfsr[95]^lfsr[101]^lfsr[103];
  assign  o_lfsr[429] = lfsr[65]^lfsr[67]^lfsr[73]^lfsr[74]^lfsr[75]^lfsr[82]^lfsr[92]^lfsr[94]^lfsr[100]^lfsr[102];
  assign  o_lfsr[430] = lfsr[64]^lfsr[66]^lfsr[72]^lfsr[73]^lfsr[74]^lfsr[81]^lfsr[91]^lfsr[93]^lfsr[99]^lfsr[101];
  assign  o_lfsr[431] = lfsr[63]^lfsr[65]^lfsr[71]^lfsr[72]^lfsr[73]^lfsr[80]^lfsr[90]^lfsr[92]^lfsr[98]^lfsr[100];
  assign  o_lfsr[432] = lfsr[62]^lfsr[64]^lfsr[70]^lfsr[71]^lfsr[72]^lfsr[79]^lfsr[89]^lfsr[91]^lfsr[97]^lfsr[99];
  assign  o_lfsr[433] = lfsr[61]^lfsr[63]^lfsr[69]^lfsr[70]^lfsr[71]^lfsr[78]^lfsr[88]^lfsr[90]^lfsr[96]^lfsr[98];
  assign  o_lfsr[434] = lfsr[60]^lfsr[62]^lfsr[68]^lfsr[69]^lfsr[70]^lfsr[77]^lfsr[87]^lfsr[89]^lfsr[95]^lfsr[97];
  assign  o_lfsr[435] = lfsr[59]^lfsr[61]^lfsr[67]^lfsr[68]^lfsr[69]^lfsr[76]^lfsr[86]^lfsr[88]^lfsr[94]^lfsr[96];
  assign  o_lfsr[436] = lfsr[58]^lfsr[60]^lfsr[66]^lfsr[67]^lfsr[68]^lfsr[75]^lfsr[85]^lfsr[87]^lfsr[93]^lfsr[95];
  assign  o_lfsr[437] = lfsr[57]^lfsr[59]^lfsr[65]^lfsr[66]^lfsr[67]^lfsr[74]^lfsr[84]^lfsr[86]^lfsr[92]^lfsr[94];
  assign  o_lfsr[438] = lfsr[56]^lfsr[58]^lfsr[64]^lfsr[65]^lfsr[66]^lfsr[73]^lfsr[83]^lfsr[85]^lfsr[91]^lfsr[93];
  assign  o_lfsr[439] = lfsr[55]^lfsr[57]^lfsr[63]^lfsr[64]^lfsr[65]^lfsr[72]^lfsr[82]^lfsr[84]^lfsr[90]^lfsr[92];
  assign  o_lfsr[440] = lfsr[54]^lfsr[56]^lfsr[62]^lfsr[63]^lfsr[64]^lfsr[71]^lfsr[81]^lfsr[83]^lfsr[89]^lfsr[91];
  assign  o_lfsr[441] = lfsr[53]^lfsr[55]^lfsr[61]^lfsr[62]^lfsr[63]^lfsr[70]^lfsr[80]^lfsr[82]^lfsr[88]^lfsr[90];
  assign  o_lfsr[442] = lfsr[52]^lfsr[54]^lfsr[60]^lfsr[61]^lfsr[62]^lfsr[69]^lfsr[79]^lfsr[81]^lfsr[87]^lfsr[89];
  assign  o_lfsr[443] = lfsr[51]^lfsr[53]^lfsr[59]^lfsr[60]^lfsr[61]^lfsr[68]^lfsr[78]^lfsr[80]^lfsr[86]^lfsr[88];
  assign  o_lfsr[444] = lfsr[50]^lfsr[52]^lfsr[58]^lfsr[59]^lfsr[60]^lfsr[67]^lfsr[77]^lfsr[79]^lfsr[85]^lfsr[87];
  assign  o_lfsr[445] = lfsr[49]^lfsr[51]^lfsr[57]^lfsr[58]^lfsr[59]^lfsr[66]^lfsr[76]^lfsr[78]^lfsr[84]^lfsr[86];
  assign  o_lfsr[446] = lfsr[48]^lfsr[50]^lfsr[56]^lfsr[57]^lfsr[58]^lfsr[65]^lfsr[75]^lfsr[77]^lfsr[83]^lfsr[85];
  assign  o_lfsr[447] = lfsr[47]^lfsr[49]^lfsr[55]^lfsr[56]^lfsr[57]^lfsr[64]^lfsr[74]^lfsr[76]^lfsr[82]^lfsr[84];
  assign  o_lfsr[448] = lfsr[46]^lfsr[48]^lfsr[54]^lfsr[55]^lfsr[56]^lfsr[63]^lfsr[73]^lfsr[75]^lfsr[81]^lfsr[83];
  assign  o_lfsr[449] = lfsr[45]^lfsr[47]^lfsr[53]^lfsr[54]^lfsr[55]^lfsr[62]^lfsr[72]^lfsr[74]^lfsr[80]^lfsr[82];
  assign  o_lfsr[450] = lfsr[44]^lfsr[46]^lfsr[52]^lfsr[53]^lfsr[54]^lfsr[61]^lfsr[71]^lfsr[73]^lfsr[79]^lfsr[81];
  assign  o_lfsr[451] = lfsr[43]^lfsr[45]^lfsr[51]^lfsr[52]^lfsr[53]^lfsr[60]^lfsr[70]^lfsr[72]^lfsr[78]^lfsr[80];
  assign  o_lfsr[452] = lfsr[42]^lfsr[44]^lfsr[50]^lfsr[51]^lfsr[52]^lfsr[59]^lfsr[69]^lfsr[71]^lfsr[77]^lfsr[79];
  assign  o_lfsr[453] = lfsr[41]^lfsr[43]^lfsr[49]^lfsr[50]^lfsr[51]^lfsr[58]^lfsr[68]^lfsr[70]^lfsr[76]^lfsr[78];
  assign  o_lfsr[454] = lfsr[40]^lfsr[42]^lfsr[48]^lfsr[49]^lfsr[50]^lfsr[57]^lfsr[67]^lfsr[69]^lfsr[75]^lfsr[77];
  assign  o_lfsr[455] = lfsr[39]^lfsr[41]^lfsr[47]^lfsr[48]^lfsr[49]^lfsr[56]^lfsr[66]^lfsr[68]^lfsr[74]^lfsr[76];
  assign  o_lfsr[456] = lfsr[38]^lfsr[40]^lfsr[46]^lfsr[47]^lfsr[48]^lfsr[55]^lfsr[65]^lfsr[67]^lfsr[73]^lfsr[75];
  assign  o_lfsr[457] = lfsr[37]^lfsr[39]^lfsr[45]^lfsr[46]^lfsr[47]^lfsr[54]^lfsr[64]^lfsr[66]^lfsr[72]^lfsr[74];
  assign  o_lfsr[458] = lfsr[36]^lfsr[38]^lfsr[44]^lfsr[45]^lfsr[46]^lfsr[53]^lfsr[63]^lfsr[65]^lfsr[71]^lfsr[73];
  assign  o_lfsr[459] = lfsr[35]^lfsr[37]^lfsr[43]^lfsr[44]^lfsr[45]^lfsr[52]^lfsr[62]^lfsr[64]^lfsr[70]^lfsr[72];
  assign  o_lfsr[460] = lfsr[34]^lfsr[36]^lfsr[42]^lfsr[43]^lfsr[44]^lfsr[51]^lfsr[61]^lfsr[63]^lfsr[69]^lfsr[71];
  assign  o_lfsr[461] = lfsr[33]^lfsr[35]^lfsr[41]^lfsr[42]^lfsr[43]^lfsr[50]^lfsr[60]^lfsr[62]^lfsr[68]^lfsr[70];
  assign  o_lfsr[462] = lfsr[32]^lfsr[34]^lfsr[40]^lfsr[41]^lfsr[42]^lfsr[49]^lfsr[59]^lfsr[61]^lfsr[67]^lfsr[69];
  assign  o_lfsr[463] = lfsr[31]^lfsr[33]^lfsr[39]^lfsr[40]^lfsr[41]^lfsr[48]^lfsr[58]^lfsr[60]^lfsr[66]^lfsr[68];
  assign  o_lfsr[464] = lfsr[30]^lfsr[32]^lfsr[38]^lfsr[39]^lfsr[40]^lfsr[47]^lfsr[57]^lfsr[59]^lfsr[65]^lfsr[67];
  assign  o_lfsr[465] = lfsr[29]^lfsr[31]^lfsr[37]^lfsr[38]^lfsr[39]^lfsr[46]^lfsr[56]^lfsr[58]^lfsr[64]^lfsr[66];
  assign  o_lfsr[466] = lfsr[28]^lfsr[30]^lfsr[36]^lfsr[37]^lfsr[38]^lfsr[45]^lfsr[55]^lfsr[57]^lfsr[63]^lfsr[65];
  assign  o_lfsr[467] = lfsr[27]^lfsr[29]^lfsr[35]^lfsr[36]^lfsr[37]^lfsr[44]^lfsr[54]^lfsr[56]^lfsr[62]^lfsr[64];
  assign  o_lfsr[468] = lfsr[26]^lfsr[28]^lfsr[34]^lfsr[35]^lfsr[36]^lfsr[43]^lfsr[53]^lfsr[55]^lfsr[61]^lfsr[63];
  assign  o_lfsr[469] = lfsr[25]^lfsr[27]^lfsr[33]^lfsr[34]^lfsr[35]^lfsr[42]^lfsr[52]^lfsr[54]^lfsr[60]^lfsr[62];
  assign  o_lfsr[470] = lfsr[24]^lfsr[26]^lfsr[32]^lfsr[33]^lfsr[34]^lfsr[41]^lfsr[51]^lfsr[53]^lfsr[59]^lfsr[61];
  assign  o_lfsr[471] = lfsr[23]^lfsr[25]^lfsr[31]^lfsr[32]^lfsr[33]^lfsr[40]^lfsr[50]^lfsr[52]^lfsr[58]^lfsr[60];
  assign  o_lfsr[472] = lfsr[22]^lfsr[24]^lfsr[30]^lfsr[31]^lfsr[32]^lfsr[39]^lfsr[49]^lfsr[51]^lfsr[57]^lfsr[59];
  assign  o_lfsr[473] = lfsr[21]^lfsr[23]^lfsr[29]^lfsr[30]^lfsr[31]^lfsr[38]^lfsr[48]^lfsr[50]^lfsr[56]^lfsr[58];
  assign  o_lfsr[474] = lfsr[20]^lfsr[22]^lfsr[28]^lfsr[29]^lfsr[30]^lfsr[37]^lfsr[47]^lfsr[49]^lfsr[55]^lfsr[57];
  assign  o_lfsr[475] = lfsr[19]^lfsr[21]^lfsr[27]^lfsr[28]^lfsr[29]^lfsr[36]^lfsr[46]^lfsr[48]^lfsr[54]^lfsr[56];
  assign  o_lfsr[476] = lfsr[18]^lfsr[20]^lfsr[26]^lfsr[27]^lfsr[28]^lfsr[35]^lfsr[45]^lfsr[47]^lfsr[53]^lfsr[55];
  assign  o_lfsr[477] = lfsr[17]^lfsr[19]^lfsr[25]^lfsr[26]^lfsr[27]^lfsr[34]^lfsr[44]^lfsr[46]^lfsr[52]^lfsr[54];
  assign  o_lfsr[478] = lfsr[16]^lfsr[18]^lfsr[24]^lfsr[25]^lfsr[26]^lfsr[33]^lfsr[43]^lfsr[45]^lfsr[51]^lfsr[53];
  assign  o_lfsr[479] = lfsr[15]^lfsr[17]^lfsr[23]^lfsr[24]^lfsr[25]^lfsr[32]^lfsr[42]^lfsr[44]^lfsr[50]^lfsr[52];
  assign  o_lfsr[480] = lfsr[14]^lfsr[16]^lfsr[22]^lfsr[23]^lfsr[24]^lfsr[31]^lfsr[41]^lfsr[43]^lfsr[49]^lfsr[51];
  assign  o_lfsr[481] = lfsr[13]^lfsr[15]^lfsr[21]^lfsr[22]^lfsr[23]^lfsr[30]^lfsr[40]^lfsr[42]^lfsr[48]^lfsr[50];
  assign  o_lfsr[482] = lfsr[12]^lfsr[14]^lfsr[20]^lfsr[21]^lfsr[22]^lfsr[29]^lfsr[39]^lfsr[41]^lfsr[47]^lfsr[49];
  assign  o_lfsr[483] = lfsr[11]^lfsr[13]^lfsr[19]^lfsr[20]^lfsr[21]^lfsr[28]^lfsr[38]^lfsr[40]^lfsr[46]^lfsr[48];
  assign  o_lfsr[484] = lfsr[10]^lfsr[12]^lfsr[18]^lfsr[19]^lfsr[20]^lfsr[27]^lfsr[37]^lfsr[39]^lfsr[45]^lfsr[47];
  assign  o_lfsr[485] = lfsr[ 9]^lfsr[11]^lfsr[17]^lfsr[18]^lfsr[19]^lfsr[26]^lfsr[36]^lfsr[38]^lfsr[44]^lfsr[46];
  assign  o_lfsr[486] = lfsr[ 8]^lfsr[10]^lfsr[16]^lfsr[17]^lfsr[18]^lfsr[25]^lfsr[35]^lfsr[37]^lfsr[43]^lfsr[45];
  assign  o_lfsr[487] = lfsr[ 7]^lfsr[ 9]^lfsr[15]^lfsr[16]^lfsr[17]^lfsr[24]^lfsr[34]^lfsr[36]^lfsr[42]^lfsr[44];
  assign  o_lfsr[488] = lfsr[ 6]^lfsr[ 8]^lfsr[14]^lfsr[15]^lfsr[16]^lfsr[23]^lfsr[33]^lfsr[35]^lfsr[41]^lfsr[43];
  assign  o_lfsr[489] = lfsr[ 5]^lfsr[ 7]^lfsr[13]^lfsr[14]^lfsr[15]^lfsr[22]^lfsr[32]^lfsr[34]^lfsr[40]^lfsr[42];
  assign  o_lfsr[490] = lfsr[ 4]^lfsr[ 6]^lfsr[12]^lfsr[13]^lfsr[14]^lfsr[21]^lfsr[31]^lfsr[33]^lfsr[39]^lfsr[41];
  assign  o_lfsr[491] = lfsr[ 3]^lfsr[ 5]^lfsr[11]^lfsr[12]^lfsr[13]^lfsr[20]^lfsr[30]^lfsr[32]^lfsr[38]^lfsr[40];
  assign  o_lfsr[492] = lfsr[ 2]^lfsr[ 4]^lfsr[10]^lfsr[11]^lfsr[12]^lfsr[19]^lfsr[29]^lfsr[31]^lfsr[37]^lfsr[39];
  assign  o_lfsr[493] = lfsr[ 1]^lfsr[ 3]^lfsr[ 9]^lfsr[10]^lfsr[11]^lfsr[18]^lfsr[28]^lfsr[30]^lfsr[36]^lfsr[38];
  assign  o_lfsr[494] = lfsr[ 0]^lfsr[ 2]^lfsr[ 8]^lfsr[ 9]^lfsr[10]^lfsr[17]^lfsr[27]^lfsr[29]^lfsr[35]^lfsr[37];
  assign  o_lfsr[495] = lfsr[ 1]^lfsr[ 7]^lfsr[ 8]^lfsr[ 9]^lfsr[16]^lfsr[26]^lfsr[28]^lfsr[34]^lfsr[36]^lfsr[98]^lfsr[100]^lfsr[125]^lfsr[127];
  assign  o_lfsr[496] = lfsr[ 0]^lfsr[ 6]^lfsr[ 7]^lfsr[ 8]^lfsr[15]^lfsr[25]^lfsr[27]^lfsr[33]^lfsr[35]^lfsr[97]^lfsr[99]^lfsr[124]^lfsr[126];
  assign  o_lfsr[497] = lfsr[ 5]^lfsr[ 6]^lfsr[ 7]^lfsr[14]^lfsr[24]^lfsr[26]^lfsr[32]^lfsr[34]^lfsr[96]^lfsr[100]^lfsr[123]^lfsr[127];
  assign  o_lfsr[498] = lfsr[ 4]^lfsr[ 5]^lfsr[ 6]^lfsr[13]^lfsr[23]^lfsr[25]^lfsr[31]^lfsr[33]^lfsr[95]^lfsr[99]^lfsr[122]^lfsr[126];
  assign  o_lfsr[499] = lfsr[ 3]^lfsr[ 4]^lfsr[ 5]^lfsr[12]^lfsr[22]^lfsr[24]^lfsr[30]^lfsr[32]^lfsr[94]^lfsr[98]^lfsr[121]^lfsr[125];
  assign  o_lfsr[500] = lfsr[ 2]^lfsr[ 3]^lfsr[ 4]^lfsr[11]^lfsr[21]^lfsr[23]^lfsr[29]^lfsr[31]^lfsr[93]^lfsr[97]^lfsr[120]^lfsr[124];
  assign  o_lfsr[501] = lfsr[ 1]^lfsr[ 2]^lfsr[ 3]^lfsr[10]^lfsr[20]^lfsr[22]^lfsr[28]^lfsr[30]^lfsr[92]^lfsr[96]^lfsr[119]^lfsr[123];
  assign  o_lfsr[502] = lfsr[ 0]^lfsr[ 1]^lfsr[ 2]^lfsr[ 9]^lfsr[19]^lfsr[21]^lfsr[27]^lfsr[29]^lfsr[91]^lfsr[95]^lfsr[118]^lfsr[122];
  assign  o_lfsr[503] = lfsr[ 0]^lfsr[ 1]^lfsr[ 8]^lfsr[18]^lfsr[20]^lfsr[26]^lfsr[28]^lfsr[90]^lfsr[94]^lfsr[98]^lfsr[100]^lfsr[117]^lfsr[121]^lfsr[125]^lfsr[127];
  assign  o_lfsr[504] = lfsr[ 0]^lfsr[ 7]^lfsr[17]^lfsr[19]^lfsr[25]^lfsr[27]^lfsr[89]^lfsr[93]^lfsr[97]^lfsr[98]^lfsr[99]^lfsr[100]^lfsr[116]^lfsr[120]^lfsr[124]^lfsr[125]^lfsr[126]^lfsr[127];
  assign  o_lfsr[505] = lfsr[ 6]^lfsr[16]^lfsr[18]^lfsr[24]^lfsr[26]^lfsr[88]^lfsr[92]^lfsr[96]^lfsr[97]^lfsr[99]^lfsr[100]^lfsr[115]^lfsr[119]^lfsr[123]^lfsr[124]^lfsr[126]^lfsr[127];
  assign  o_lfsr[506] = lfsr[ 5]^lfsr[15]^lfsr[17]^lfsr[23]^lfsr[25]^lfsr[87]^lfsr[91]^lfsr[95]^lfsr[96]^lfsr[98]^lfsr[99]^lfsr[114]^lfsr[118]^lfsr[122]^lfsr[123]^lfsr[125]^lfsr[126];
  assign  o_lfsr[507] = lfsr[ 4]^lfsr[14]^lfsr[16]^lfsr[22]^lfsr[24]^lfsr[86]^lfsr[90]^lfsr[94]^lfsr[95]^lfsr[97]^lfsr[98]^lfsr[113]^lfsr[117]^lfsr[121]^lfsr[122]^lfsr[124]^lfsr[125];
  assign  o_lfsr[508] = lfsr[ 3]^lfsr[13]^lfsr[15]^lfsr[21]^lfsr[23]^lfsr[85]^lfsr[89]^lfsr[93]^lfsr[94]^lfsr[96]^lfsr[97]^lfsr[112]^lfsr[116]^lfsr[120]^lfsr[121]^lfsr[123]^lfsr[124];
  assign  o_lfsr[509] = lfsr[ 2]^lfsr[12]^lfsr[14]^lfsr[20]^lfsr[22]^lfsr[84]^lfsr[88]^lfsr[92]^lfsr[93]^lfsr[95]^lfsr[96]^lfsr[111]^lfsr[115]^lfsr[119]^lfsr[120]^lfsr[122]^lfsr[123];
  assign  o_lfsr[510] = lfsr[ 1]^lfsr[11]^lfsr[13]^lfsr[19]^lfsr[21]^lfsr[83]^lfsr[87]^lfsr[91]^lfsr[92]^lfsr[94]^lfsr[95]^lfsr[110]^lfsr[114]^lfsr[118]^lfsr[119]^lfsr[121]^lfsr[122];
  assign  o_lfsr[511] = lfsr[ 0]^lfsr[10]^lfsr[12]^lfsr[18]^lfsr[20]^lfsr[82]^lfsr[86]^lfsr[90]^lfsr[91]^lfsr[93]^lfsr[94]^lfsr[109]^lfsr[113]^lfsr[117]^lfsr[118]^lfsr[120]^lfsr[121];

  // To advance the state by N=512 clocks:
  localparam N=512;

  always @(posedge(clk)) begin : lfsr_clock
    if (reset == 1'b1) begin
       lfsr <= {(512){1'b1}};
    end else begin
       if (i_init==1'b1) begin
          lfsr <= i_seed;
       end else begin
          if (i_advance==1'b1) begin
             for (i=0; i<128; i=i+1) begin
                lfsr[i]  <= (N-1>=i) ? o_lfsr[N-1-i]:lfsr[i-N];
             end
          end
       end
    end
  end // always

endmodule  // lfsr

`default_nettype wire

